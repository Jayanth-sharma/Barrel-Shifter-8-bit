magic
tech scmos
magscale 1 2
timestamp 1668920897
<< metal1 >>
rect 248 806 254 814
rect 262 806 268 814
rect 276 806 282 814
rect 290 806 296 814
rect 164 716 172 724
rect 189 703 195 723
rect 29 697 67 703
rect 125 697 163 703
rect 189 697 227 703
rect 429 703 435 723
rect 244 697 307 703
rect 349 697 403 703
rect 429 697 467 703
rect 509 697 547 703
rect 605 697 643 703
rect 653 697 691 703
rect 845 697 883 703
rect 989 697 1004 703
rect 237 677 284 683
rect 484 677 499 683
rect 93 657 115 663
rect 493 657 499 677
rect 573 677 588 683
rect 909 677 924 683
rect 964 677 979 683
rect 973 657 979 677
rect 804 636 806 644
rect 728 606 734 614
rect 742 606 748 614
rect 756 606 762 614
rect 770 606 776 614
rect 36 576 38 584
rect 874 576 876 584
rect 141 543 147 556
rect 125 537 147 543
rect 324 537 339 543
rect 477 537 483 563
rect 573 537 588 543
rect 845 537 860 543
rect 157 517 195 523
rect 221 517 259 523
rect 45 497 60 503
rect 221 497 227 517
rect 308 517 355 523
rect 381 517 419 523
rect 381 497 387 517
rect 573 517 611 523
rect 733 517 780 523
rect 461 497 476 503
rect 573 497 579 517
rect 1012 517 1027 523
rect 826 436 828 444
rect 248 406 254 414
rect 262 406 268 414
rect 276 406 282 414
rect 290 406 296 414
rect 404 376 406 384
rect 77 297 115 303
rect 125 297 163 303
rect 429 303 435 323
rect 365 297 403 303
rect 429 297 444 303
rect 621 303 627 323
rect 557 297 595 303
rect 621 297 659 303
rect 797 297 835 303
rect 221 277 268 283
rect 621 277 636 283
rect 333 257 355 263
rect 458 236 460 244
rect 708 236 710 244
rect 728 206 734 214
rect 742 206 748 214
rect 756 206 762 214
rect 770 206 776 214
rect 93 157 115 163
rect 301 144 307 163
rect 237 137 300 143
rect 573 137 595 143
rect 29 117 67 123
rect 125 117 163 123
rect 509 117 547 123
rect 813 117 851 123
rect 868 117 883 123
rect 1012 117 1027 123
rect 248 6 254 14
rect 262 6 268 14
rect 276 6 282 14
rect 290 6 296 14
<< m2contact >>
rect 254 806 262 814
rect 268 806 276 814
rect 282 806 290 814
rect 332 776 340 784
rect 716 776 724 784
rect 92 716 100 724
rect 156 716 164 724
rect 204 716 212 724
rect 236 696 244 704
rect 444 716 452 724
rect 572 716 580 724
rect 668 716 676 724
rect 812 716 820 724
rect 908 716 916 724
rect 924 716 932 724
rect 1004 716 1012 724
rect 1004 696 1012 704
rect 1036 696 1044 704
rect 44 676 52 684
rect 140 676 148 684
rect 284 676 292 684
rect 380 676 388 684
rect 412 676 420 684
rect 476 676 484 684
rect 12 656 20 664
rect 364 656 372 664
rect 524 676 532 684
rect 588 676 596 684
rect 620 676 628 684
rect 780 676 788 684
rect 860 676 868 684
rect 924 676 932 684
rect 956 676 964 684
rect 588 656 596 664
rect 828 656 836 664
rect 1020 676 1028 684
rect 1052 676 1060 684
rect 796 636 804 644
rect 924 636 932 644
rect 734 606 742 614
rect 748 606 756 614
rect 762 606 770 614
rect 28 576 36 584
rect 220 576 228 584
rect 428 576 436 584
rect 508 576 516 584
rect 668 576 676 584
rect 876 576 884 584
rect 892 576 900 584
rect 908 576 916 584
rect 940 576 948 584
rect 60 556 68 564
rect 140 556 148 564
rect 380 556 388 564
rect 444 556 452 564
rect 12 536 20 544
rect 172 536 180 544
rect 268 536 276 544
rect 316 536 324 544
rect 428 536 436 544
rect 684 556 692 564
rect 716 556 724 564
rect 524 536 532 544
rect 588 536 596 544
rect 620 536 628 544
rect 636 536 644 544
rect 860 536 868 544
rect 892 536 900 544
rect 908 536 916 544
rect 1004 536 1012 544
rect 60 496 68 504
rect 76 496 84 504
rect 92 496 100 504
rect 300 516 308 524
rect 236 496 244 504
rect 540 516 548 524
rect 396 496 404 504
rect 476 496 484 504
rect 508 496 516 504
rect 780 516 788 524
rect 828 516 836 524
rect 972 516 980 524
rect 988 516 996 524
rect 1004 516 1012 524
rect 588 496 596 504
rect 668 496 676 504
rect 700 496 708 504
rect 796 496 804 504
rect 860 496 868 504
rect 940 496 948 504
rect 956 496 964 504
rect 1052 476 1060 484
rect 108 436 116 444
rect 828 436 836 444
rect 254 406 262 414
rect 268 406 276 414
rect 282 406 290 414
rect 396 376 404 384
rect 940 376 948 384
rect 44 336 52 344
rect 1052 336 1060 344
rect 92 316 100 324
rect 188 316 196 324
rect 332 316 340 324
rect 28 296 36 304
rect 300 296 308 304
rect 444 316 452 324
rect 524 316 532 324
rect 444 296 452 304
rect 636 316 644 324
rect 716 316 724 324
rect 860 316 868 324
rect 908 316 916 324
rect 956 316 964 324
rect 972 296 980 304
rect 1020 296 1028 304
rect 140 276 148 284
rect 268 276 276 284
rect 284 276 292 284
rect 316 276 324 284
rect 380 276 388 284
rect 476 276 484 284
rect 492 276 500 284
rect 572 276 580 284
rect 636 276 644 284
rect 668 276 676 284
rect 684 276 692 284
rect 812 276 820 284
rect 860 276 868 284
rect 876 276 884 284
rect 924 276 932 284
rect 1004 276 1012 284
rect 12 256 20 264
rect 172 256 180 264
rect 508 256 516 264
rect 540 256 548 264
rect 780 256 788 264
rect 188 236 196 244
rect 460 236 468 244
rect 476 236 484 244
rect 492 236 500 244
rect 668 236 676 244
rect 700 236 708 244
rect 908 236 916 244
rect 734 206 742 214
rect 748 206 756 214
rect 762 206 770 214
rect 332 176 340 184
rect 444 176 452 184
rect 12 156 20 164
rect 428 156 436 164
rect 492 156 500 164
rect 636 156 644 164
rect 860 156 868 164
rect 924 156 932 164
rect 44 136 52 144
rect 140 136 148 144
rect 172 136 180 144
rect 300 136 308 144
rect 364 136 372 144
rect 380 136 388 144
rect 476 136 484 144
rect 524 136 532 144
rect 556 136 564 144
rect 684 136 692 144
rect 716 136 724 144
rect 828 136 836 144
rect 1004 136 1012 144
rect 316 116 324 124
rect 396 116 404 124
rect 700 116 708 124
rect 796 116 804 124
rect 860 116 868 124
rect 972 116 980 124
rect 988 116 996 124
rect 1004 116 1012 124
rect 92 96 100 104
rect 188 96 196 104
rect 204 96 212 104
rect 220 96 228 104
rect 332 96 340 104
rect 428 96 436 104
rect 444 96 452 104
rect 572 96 580 104
rect 620 96 628 104
rect 652 96 660 104
rect 668 96 676 104
rect 780 96 788 104
rect 940 96 948 104
rect 956 96 964 104
rect 604 76 612 84
rect 1052 76 1060 84
rect 908 36 916 44
rect 254 6 262 14
rect 268 6 276 14
rect 282 6 290 14
<< metal2 >>
rect 301 837 339 843
rect 349 837 371 843
rect 248 806 254 814
rect 262 806 268 814
rect 276 806 282 814
rect 290 806 296 814
rect 333 784 339 837
rect 13 664 19 696
rect 29 584 35 716
rect 13 544 19 556
rect 45 524 51 676
rect 157 583 163 716
rect 205 684 211 716
rect 141 577 163 583
rect 141 564 147 577
rect 61 504 67 516
rect 93 504 99 536
rect 45 324 51 336
rect 13 264 19 276
rect 13 104 19 156
rect 61 144 67 496
rect 109 323 115 436
rect 100 317 115 323
rect 141 284 147 536
rect 189 264 195 316
rect 205 264 211 676
rect 237 583 243 696
rect 365 664 371 837
rect 397 683 403 716
rect 445 684 451 716
rect 477 684 483 843
rect 701 837 723 843
rect 717 784 723 837
rect 781 804 787 843
rect 813 724 819 796
rect 388 677 403 683
rect 228 577 243 583
rect 269 544 275 656
rect 237 524 243 536
rect 237 504 243 516
rect 269 444 275 536
rect 301 504 307 516
rect 317 504 323 536
rect 397 504 403 677
rect 413 584 419 676
rect 509 584 515 716
rect 605 677 620 683
rect 429 544 435 576
rect 445 564 451 576
rect 248 406 254 414
rect 262 406 268 414
rect 276 406 282 414
rect 290 406 296 414
rect 317 324 323 496
rect 397 384 403 436
rect 509 324 515 496
rect 525 484 531 536
rect 605 524 611 677
rect 669 584 675 716
rect 813 684 819 716
rect 728 606 734 614
rect 742 606 748 614
rect 756 606 762 614
rect 770 606 776 614
rect 621 544 627 556
rect 717 544 723 556
rect 541 504 547 516
rect 669 504 675 516
rect 589 484 595 496
rect 589 324 595 476
rect 717 324 723 516
rect 797 504 803 636
rect 861 544 867 676
rect 877 584 883 716
rect 893 544 899 576
rect 909 544 915 576
rect 829 504 835 516
rect 861 504 867 536
rect 861 484 867 496
rect 829 344 835 436
rect 285 284 291 316
rect 141 144 147 256
rect 173 144 179 256
rect 189 104 195 236
rect 333 184 339 316
rect 381 264 387 276
rect 445 184 451 296
rect 477 244 483 276
rect 493 244 499 276
rect 509 244 515 256
rect 365 144 371 176
rect 205 104 211 136
rect 301 43 307 136
rect 333 104 339 136
rect 301 37 323 43
rect 248 6 254 14
rect 262 6 268 14
rect 276 6 282 14
rect 290 6 296 14
rect 317 -17 323 37
rect 365 -17 371 136
rect 445 104 451 116
rect 461 104 467 236
rect 493 164 499 176
rect 477 144 483 156
rect 525 144 531 316
rect 573 284 579 316
rect 717 304 723 316
rect 813 284 819 296
rect 573 264 579 276
rect 548 257 563 263
rect 557 144 563 257
rect 573 104 579 236
rect 621 124 627 256
rect 669 244 675 276
rect 781 264 787 276
rect 685 144 691 156
rect 701 144 707 236
rect 728 206 734 214
rect 742 206 748 214
rect 756 206 762 214
rect 770 206 776 214
rect 829 144 835 296
rect 877 284 883 336
rect 925 324 931 636
rect 941 584 947 736
rect 1005 724 1011 736
rect 1053 684 1059 716
rect 1005 544 1011 676
rect 941 504 947 536
rect 989 504 995 516
rect 941 463 947 496
rect 957 484 963 496
rect 941 457 963 463
rect 941 384 947 436
rect 957 324 963 457
rect 909 304 915 316
rect 957 304 963 316
rect 1021 304 1027 676
rect 1053 484 1059 496
rect 877 163 883 276
rect 868 157 883 163
rect 717 124 723 136
rect 621 104 627 116
rect 701 104 707 116
rect 781 104 787 136
rect 909 124 915 236
rect 925 164 931 276
rect 957 144 963 296
rect 973 284 979 296
rect 1005 284 1011 296
rect 957 104 963 116
rect 989 104 995 116
rect 669 84 675 96
rect 1053 84 1059 96
rect 909 -17 915 36
rect 301 -23 323 -17
rect 349 -23 371 -17
rect 893 -23 915 -17
<< m3contact >>
rect 254 806 262 814
rect 268 806 276 814
rect 282 806 290 814
rect 28 716 36 724
rect 92 716 100 724
rect 12 696 20 704
rect 140 676 148 684
rect 12 556 20 564
rect 204 676 212 684
rect 60 556 68 564
rect 92 536 100 544
rect 140 536 148 544
rect 172 536 180 544
rect 44 516 52 524
rect 60 516 68 524
rect 76 496 84 504
rect 44 316 52 324
rect 28 296 36 304
rect 12 276 20 284
rect 284 676 292 684
rect 396 716 404 724
rect 444 716 452 724
rect 780 796 788 804
rect 812 796 820 804
rect 940 736 948 744
rect 1004 736 1012 744
rect 508 716 516 724
rect 572 716 580 724
rect 876 716 884 724
rect 908 716 916 724
rect 924 716 932 724
rect 268 656 276 664
rect 380 556 388 564
rect 236 536 244 544
rect 236 516 244 524
rect 412 676 420 684
rect 444 676 452 684
rect 524 676 532 684
rect 588 676 596 684
rect 588 656 596 664
rect 412 576 420 584
rect 444 576 452 584
rect 588 536 596 544
rect 300 496 308 504
rect 316 496 324 504
rect 396 496 404 504
rect 476 496 484 504
rect 268 436 276 444
rect 254 406 262 414
rect 268 406 276 414
rect 282 406 290 414
rect 396 436 404 444
rect 780 676 788 684
rect 812 676 820 684
rect 860 676 868 684
rect 828 656 836 664
rect 734 606 742 614
rect 748 606 756 614
rect 762 606 770 614
rect 620 556 628 564
rect 684 556 692 564
rect 636 536 644 544
rect 716 536 724 544
rect 604 516 612 524
rect 668 516 676 524
rect 716 516 724 524
rect 780 516 788 524
rect 540 496 548 504
rect 700 496 708 504
rect 524 476 532 484
rect 588 476 596 484
rect 924 676 932 684
rect 828 496 836 504
rect 860 476 868 484
rect 828 336 836 344
rect 876 336 884 344
rect 284 316 292 324
rect 316 316 324 324
rect 444 316 452 324
rect 508 316 516 324
rect 524 316 532 324
rect 572 316 580 324
rect 588 316 596 324
rect 636 316 644 324
rect 860 316 868 324
rect 300 296 308 304
rect 268 276 276 284
rect 316 276 324 284
rect 140 256 148 264
rect 188 256 196 264
rect 204 256 212 264
rect 44 136 52 144
rect 60 136 68 144
rect 380 256 388 264
rect 508 236 516 244
rect 364 176 372 184
rect 428 156 436 164
rect 204 136 212 144
rect 332 136 340 144
rect 380 136 388 144
rect 12 96 20 104
rect 92 96 100 104
rect 220 96 228 104
rect 316 116 324 124
rect 254 6 262 14
rect 268 6 276 14
rect 282 6 290 14
rect 396 116 404 124
rect 444 116 452 124
rect 492 176 500 184
rect 476 156 484 164
rect 716 296 724 304
rect 812 296 820 304
rect 828 296 836 304
rect 636 276 644 284
rect 684 276 692 284
rect 780 276 788 284
rect 572 256 580 264
rect 620 256 628 264
rect 572 236 580 244
rect 524 136 532 144
rect 636 156 644 164
rect 684 156 692 164
rect 734 206 742 214
rect 748 206 756 214
rect 762 206 770 214
rect 1052 716 1060 724
rect 1004 696 1012 704
rect 1036 696 1044 704
rect 956 676 964 684
rect 1004 676 1012 684
rect 1052 676 1060 684
rect 940 536 948 544
rect 1004 536 1012 544
rect 972 516 980 524
rect 1004 516 1012 524
rect 988 496 996 504
rect 956 476 964 484
rect 940 436 948 444
rect 924 316 932 324
rect 1052 496 1060 504
rect 1052 336 1060 344
rect 908 296 916 304
rect 956 296 964 304
rect 1004 296 1012 304
rect 860 276 868 284
rect 700 136 708 144
rect 780 136 788 144
rect 620 116 628 124
rect 716 116 724 124
rect 924 156 932 164
rect 972 276 980 284
rect 956 136 964 144
rect 1004 136 1012 144
rect 796 116 804 124
rect 860 116 868 124
rect 908 116 916 124
rect 956 116 964 124
rect 972 116 980 124
rect 1004 116 1012 124
rect 428 96 436 104
rect 460 96 468 104
rect 652 96 660 104
rect 700 96 708 104
rect 940 96 948 104
rect 988 96 996 104
rect 1052 96 1060 104
rect 604 76 612 84
rect 668 76 676 84
<< metal3 >>
rect 248 814 296 816
rect 248 806 252 814
rect 262 806 268 814
rect 276 806 282 814
rect 292 806 296 814
rect 248 804 296 806
rect 788 797 812 803
rect 948 737 1004 743
rect 36 717 92 723
rect 404 717 444 723
rect 516 717 572 723
rect 884 717 908 723
rect 932 717 1052 723
rect -19 697 12 703
rect 1012 697 1036 703
rect 148 677 204 683
rect 292 677 412 683
rect 452 677 524 683
rect 596 677 780 683
rect 820 677 860 683
rect 932 677 956 683
rect 1012 677 1052 683
rect 1060 677 1091 683
rect 276 657 588 663
rect 781 663 787 676
rect 781 657 828 663
rect 728 614 776 616
rect 728 606 732 614
rect 742 606 748 614
rect 756 606 762 614
rect 772 606 776 614
rect 728 604 776 606
rect 420 577 444 583
rect -19 557 12 563
rect 20 557 60 563
rect 388 557 620 563
rect 628 557 684 563
rect 100 537 140 543
rect 148 537 172 543
rect 180 537 236 543
rect 596 537 636 543
rect 644 537 716 543
rect 948 537 1004 543
rect -19 517 44 523
rect 52 517 60 523
rect 244 517 604 523
rect 612 517 668 523
rect 676 517 716 523
rect 788 517 963 523
rect 84 497 300 503
rect 324 497 396 503
rect 484 497 540 503
rect 708 497 828 503
rect 957 503 963 517
rect 980 517 1004 523
rect 957 497 988 503
rect 1060 497 1091 503
rect 532 477 588 483
rect 596 477 860 483
rect 948 477 956 483
rect 276 437 396 443
rect 248 414 296 416
rect 248 406 252 414
rect 262 406 268 414
rect 276 406 282 414
rect 292 406 296 414
rect 248 404 296 406
rect 836 337 876 343
rect 1060 337 1091 343
rect -19 317 44 323
rect 292 317 316 323
rect 324 317 444 323
rect 452 317 508 323
rect 516 317 524 323
rect 580 317 588 323
rect 596 317 636 323
rect 868 317 924 323
rect 36 297 300 303
rect 724 297 812 303
rect 820 297 828 303
rect 836 297 908 303
rect 916 297 956 303
rect 1012 297 1091 303
rect -19 277 12 283
rect 276 277 316 283
rect 644 277 684 283
rect 692 277 780 283
rect 868 277 972 283
rect 148 257 188 263
rect 196 257 204 263
rect 212 257 380 263
rect 388 257 572 263
rect 580 257 620 263
rect 516 237 572 243
rect 728 214 776 216
rect 728 206 732 214
rect 742 206 748 214
rect 756 206 762 214
rect 772 206 776 214
rect 728 204 776 206
rect 372 177 492 183
rect 436 157 476 163
rect 484 157 636 163
rect 692 157 924 163
rect 52 137 60 143
rect 68 137 204 143
rect 212 137 332 143
rect 340 137 380 143
rect 388 137 524 143
rect 708 137 780 143
rect 964 137 1004 143
rect 324 117 396 123
rect 452 117 620 123
rect 628 117 716 123
rect 804 117 860 123
rect 916 117 956 123
rect 980 117 1004 123
rect -19 97 12 103
rect 100 97 220 103
rect 436 97 460 103
rect 660 97 700 103
rect 948 97 988 103
rect 1060 97 1091 103
rect 612 77 668 83
rect 248 14 296 16
rect 248 6 252 14
rect 262 6 268 14
rect 276 6 282 14
rect 292 6 296 14
rect 248 4 296 6
<< m4contact >>
rect 252 806 254 814
rect 254 806 260 814
rect 268 806 276 814
rect 284 806 290 814
rect 290 806 292 814
rect 732 606 734 614
rect 734 606 740 614
rect 748 606 756 614
rect 764 606 770 614
rect 770 606 772 614
rect 940 476 948 484
rect 940 436 948 444
rect 252 406 254 414
rect 254 406 260 414
rect 268 406 276 414
rect 284 406 290 414
rect 290 406 292 414
rect 732 206 734 214
rect 734 206 740 214
rect 748 206 756 214
rect 764 206 770 214
rect 770 206 772 214
rect 252 6 254 14
rect 254 6 260 14
rect 268 6 276 14
rect 284 6 290 14
rect 290 6 292 14
<< metal4 >>
rect 248 814 296 840
rect 248 806 252 814
rect 260 806 268 814
rect 276 806 284 814
rect 292 806 296 814
rect 248 414 296 806
rect 248 406 252 414
rect 260 406 268 414
rect 276 406 284 414
rect 292 406 296 414
rect 248 14 296 406
rect 248 6 252 14
rect 260 6 268 14
rect 276 6 284 14
rect 292 6 296 14
rect 248 -40 296 6
rect 728 614 776 840
rect 728 606 732 614
rect 740 606 748 614
rect 756 606 764 614
rect 772 606 776 614
rect 728 214 776 606
rect 938 484 950 486
rect 938 476 940 484
rect 948 476 950 484
rect 938 444 950 476
rect 938 436 940 444
rect 948 436 950 444
rect 938 434 950 436
rect 728 206 732 214
rect 740 206 748 214
rect 756 206 764 214
rect 772 206 776 214
rect 728 -40 776 206
use INVX1  INVX1_18
timestamp 1668920897
transform 1 0 8 0 -1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_19
timestamp 1668920897
transform 1 0 40 0 -1 210
box -4 -6 68 206
use INVX1  INVX1_20
timestamp 1668920897
transform 1 0 8 0 1 210
box -4 -6 36 206
use BUFX2  BUFX2_1
timestamp 1668920897
transform -1 0 88 0 1 210
box -4 -6 52 206
use INVX1  INVX1_2
timestamp 1668920897
transform 1 0 104 0 -1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_3
timestamp 1668920897
transform 1 0 136 0 -1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_11
timestamp 1668920897
transform -1 0 152 0 1 210
box -4 -6 68 206
use INVX1  INVX1_10
timestamp 1668920897
transform -1 0 184 0 1 210
box -4 -6 36 206
use NAND2X1  NAND2X1_18
timestamp 1668920897
transform -1 0 248 0 -1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_2
timestamp 1668920897
transform -1 0 232 0 1 210
box -4 -6 52 206
use FILL  FILL_0_0_0
timestamp 1668920897
transform 1 0 248 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_1
timestamp 1668920897
transform 1 0 264 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_2
timestamp 1668920897
transform 1 0 280 0 -1 210
box -4 -6 20 206
use INVX1  INVX1_22
timestamp 1668920897
transform 1 0 296 0 -1 210
box -4 -6 36 206
use FILL  FILL_1_0_0
timestamp 1668920897
transform 1 0 232 0 1 210
box -4 -6 20 206
use FILL  FILL_1_0_1
timestamp 1668920897
transform 1 0 248 0 1 210
box -4 -6 20 206
use FILL  FILL_1_0_2
timestamp 1668920897
transform 1 0 264 0 1 210
box -4 -6 20 206
use OAI21X1  OAI21X1_21
timestamp 1668920897
transform 1 0 280 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_20
timestamp 1668920897
transform -1 0 376 0 -1 210
box -4 -6 52 206
use INVX1  INVX1_4
timestamp 1668920897
transform 1 0 344 0 1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_23
timestamp 1668920897
transform 1 0 376 0 -1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_4
timestamp 1668920897
transform -1 0 488 0 -1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_5
timestamp 1668920897
transform 1 0 376 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_22
timestamp 1668920897
transform -1 0 488 0 1 210
box -4 -6 52 206
use INVX1  INVX1_24
timestamp 1668920897
transform 1 0 488 0 -1 210
box -4 -6 36 206
use NAND2X1  NAND2X1_24
timestamp 1668920897
transform 1 0 488 0 1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_1
timestamp 1668920897
transform 1 0 520 0 -1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_6
timestamp 1668920897
transform 1 0 584 0 -1 210
box -4 -6 52 206
use INVX1  INVX1_8
timestamp 1668920897
transform 1 0 536 0 1 210
box -4 -6 36 206
use OAI21X1  OAI21X1_9
timestamp 1668920897
transform 1 0 568 0 1 210
box -4 -6 68 206
use INVX1  INVX1_6
timestamp 1668920897
transform 1 0 632 0 -1 210
box -4 -6 36 206
use NAND2X1  NAND2X1_8
timestamp 1668920897
transform -1 0 680 0 1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_7
timestamp 1668920897
transform -1 0 728 0 -1 210
box -4 -6 68 206
use FILL  FILL_0_1_0
timestamp 1668920897
transform -1 0 744 0 -1 210
box -4 -6 20 206
use NAND2X1  NAND2X1_15
timestamp 1668920897
transform 1 0 680 0 1 210
box -4 -6 52 206
use FILL  FILL_1_1_0
timestamp 1668920897
transform 1 0 728 0 1 210
box -4 -6 20 206
use FILL  FILL_0_1_1
timestamp 1668920897
transform -1 0 760 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_2
timestamp 1668920897
transform -1 0 776 0 -1 210
box -4 -6 20 206
use OAI21X1  OAI21X1_16
timestamp 1668920897
transform -1 0 840 0 -1 210
box -4 -6 68 206
use FILL  FILL_1_1_1
timestamp 1668920897
transform 1 0 744 0 1 210
box -4 -6 20 206
use FILL  FILL_1_1_2
timestamp 1668920897
transform 1 0 760 0 1 210
box -4 -6 20 206
use INVX1  INVX1_16
timestamp 1668920897
transform 1 0 776 0 1 210
box -4 -6 36 206
use INVX1  INVX1_15
timestamp 1668920897
transform -1 0 872 0 -1 210
box -4 -6 36 206
use BUFX2  BUFX2_6
timestamp 1668920897
transform 1 0 872 0 -1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_17
timestamp 1668920897
transform 1 0 808 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_14
timestamp 1668920897
transform 1 0 872 0 1 210
box -4 -6 52 206
use INVX1  INVX1_14
timestamp 1668920897
transform 1 0 920 0 -1 210
box -4 -6 36 206
use NAND2X1  NAND2X1_13
timestamp 1668920897
transform 1 0 920 0 1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_15
timestamp 1668920897
transform -1 0 1016 0 -1 210
box -4 -6 68 206
use BUFX2  BUFX2_5
timestamp 1668920897
transform 1 0 1016 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_7
timestamp 1668920897
transform 1 0 968 0 1 210
box -4 -6 52 206
use BUFX2  BUFX2_8
timestamp 1668920897
transform 1 0 1016 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_19
timestamp 1668920897
transform 1 0 8 0 -1 610
box -4 -6 52 206
use INVX1  INVX1_23
timestamp 1668920897
transform 1 0 56 0 -1 610
box -4 -6 36 206
use NAND2X1  NAND2X1_10
timestamp 1668920897
transform -1 0 136 0 -1 610
box -4 -6 52 206
use INVX1  INVX1_11
timestamp 1668920897
transform 1 0 136 0 -1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_12
timestamp 1668920897
transform 1 0 168 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_11
timestamp 1668920897
transform -1 0 280 0 -1 610
box -4 -6 52 206
use FILL  FILL_2_0_0
timestamp 1668920897
transform 1 0 280 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_1
timestamp 1668920897
transform 1 0 296 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_2
timestamp 1668920897
transform 1 0 312 0 -1 610
box -4 -6 20 206
use OAI21X1  OAI21X1_24
timestamp 1668920897
transform 1 0 328 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_23
timestamp 1668920897
transform -1 0 440 0 -1 610
box -4 -6 52 206
use INVX1  INVX1_5
timestamp 1668920897
transform 1 0 440 0 -1 610
box -4 -6 36 206
use NAND2X1  NAND2X1_1
timestamp 1668920897
transform 1 0 472 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_6
timestamp 1668920897
transform 1 0 520 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_5
timestamp 1668920897
transform -1 0 632 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_12
timestamp 1668920897
transform 1 0 632 0 -1 610
box -4 -6 52 206
use INVX1  INVX1_7
timestamp 1668920897
transform 1 0 680 0 -1 610
box -4 -6 36 206
use INVX1  INVX1_13
timestamp 1668920897
transform 1 0 712 0 -1 610
box -4 -6 36 206
use FILL  FILL_2_1_0
timestamp 1668920897
transform -1 0 760 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_1
timestamp 1668920897
transform -1 0 776 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_2
timestamp 1668920897
transform -1 0 792 0 -1 610
box -4 -6 20 206
use OAI21X1  OAI21X1_8
timestamp 1668920897
transform -1 0 856 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_9
timestamp 1668920897
transform -1 0 904 0 -1 610
box -4 -6 52 206
use NAND2X1  NAND2X1_17
timestamp 1668920897
transform 1 0 904 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_14
timestamp 1668920897
transform -1 0 1016 0 -1 610
box -4 -6 68 206
use BUFX2  BUFX2_4
timestamp 1668920897
transform 1 0 1016 0 -1 610
box -4 -6 52 206
use INVX1  INVX1_19
timestamp 1668920897
transform 1 0 8 0 1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_20
timestamp 1668920897
transform 1 0 40 0 1 610
box -4 -6 68 206
use INVX1  INVX1_3
timestamp 1668920897
transform 1 0 104 0 1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_4
timestamp 1668920897
transform 1 0 136 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_3
timestamp 1668920897
transform -1 0 248 0 1 610
box -4 -6 52 206
use FILL  FILL_3_0_0
timestamp 1668920897
transform 1 0 248 0 1 610
box -4 -6 20 206
use FILL  FILL_3_0_1
timestamp 1668920897
transform 1 0 264 0 1 610
box -4 -6 20 206
use FILL  FILL_3_0_2
timestamp 1668920897
transform 1 0 280 0 1 610
box -4 -6 20 206
use BUFX2  BUFX2_2
timestamp 1668920897
transform 1 0 296 0 1 610
box -4 -6 52 206
use INVX1  INVX1_21
timestamp 1668920897
transform -1 0 376 0 1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_22
timestamp 1668920897
transform 1 0 376 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_21
timestamp 1668920897
transform -1 0 488 0 1 610
box -4 -6 52 206
use INVX1  INVX1_1
timestamp 1668920897
transform 1 0 488 0 1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_2
timestamp 1668920897
transform 1 0 520 0 1 610
box -4 -6 68 206
use INVX1  INVX1_12
timestamp 1668920897
transform 1 0 584 0 1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_13
timestamp 1668920897
transform 1 0 616 0 1 610
box -4 -6 68 206
use BUFX2  BUFX2_3
timestamp 1668920897
transform 1 0 680 0 1 610
box -4 -6 52 206
use FILL  FILL_3_1_0
timestamp 1668920897
transform 1 0 728 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1_1
timestamp 1668920897
transform 1 0 744 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1_2
timestamp 1668920897
transform 1 0 760 0 1 610
box -4 -6 20 206
use NAND2X1  NAND2X1_7
timestamp 1668920897
transform 1 0 776 0 1 610
box -4 -6 52 206
use INVX1  INVX1_9
timestamp 1668920897
transform 1 0 824 0 1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_10
timestamp 1668920897
transform 1 0 856 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_16
timestamp 1668920897
transform -1 0 968 0 1 610
box -4 -6 52 206
use INVX1  INVX1_17
timestamp 1668920897
transform 1 0 968 0 1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_18
timestamp 1668920897
transform -1 0 1064 0 1 610
box -4 -6 68 206
<< labels >>
flabel metal4 s 248 -40 296 -16 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal4 s 728 -40 776 -16 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal3 s -19 97 -13 103 7 FreeSans 24 0 0 0 in[0]
port 2 nsew
flabel metal3 s -19 697 -13 703 7 FreeSans 24 0 0 0 in[1]
port 3 nsew
flabel metal3 s -19 277 -13 283 7 FreeSans 24 0 0 0 in[2]
port 4 nsew
flabel metal2 s 349 837 355 843 3 FreeSans 24 90 0 0 in[3]
port 5 nsew
flabel metal2 s 301 -23 307 -17 7 FreeSans 24 270 0 0 in[4]
port 6 nsew
flabel metal3 s -19 557 -13 563 7 FreeSans 24 0 0 0 in[5]
port 7 nsew
flabel metal2 s 349 -23 355 -17 7 FreeSans 24 270 0 0 in[6]
port 8 nsew
flabel metal2 s 477 837 483 843 3 FreeSans 24 90 0 0 in[7]
port 9 nsew
flabel metal3 s 1085 677 1091 683 3 FreeSans 24 0 0 0 ctrl[0]
port 10 nsew
flabel metal2 s 781 837 787 843 3 FreeSans 24 90 0 0 ctrl[1]
port 11 nsew
flabel metal3 s -19 517 -13 523 7 FreeSans 24 0 0 0 ctrl[2]
port 12 nsew
flabel metal3 s -19 317 -13 323 7 FreeSans 24 0 0 0 out[0]
port 13 nsew
flabel metal2 s 301 837 307 843 3 FreeSans 24 90 0 0 out[1]
port 14 nsew
flabel metal2 s 701 837 707 843 3 FreeSans 24 90 0 0 out[2]
port 15 nsew
flabel metal3 s 1085 497 1091 503 3 FreeSans 24 0 0 0 out[3]
port 16 nsew
flabel metal3 s 1085 97 1091 103 3 FreeSans 24 0 0 0 out[4]
port 17 nsew
flabel metal2 s 893 -23 899 -17 7 FreeSans 24 270 0 0 out[5]
port 18 nsew
flabel metal3 s 1085 297 1091 303 3 FreeSans 24 0 0 0 out[6]
port 19 nsew
flabel metal3 s 1085 337 1091 343 3 FreeSans 24 0 0 0 out[7]
port 20 nsew
<< end >>
