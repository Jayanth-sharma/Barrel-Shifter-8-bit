* NGSPICE file created from barrel_shifter_8bit.ext - technology: scmos

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

.subckt barrel_shifter_8bit vdd gnd in[0] in[1] in[2] in[3] in[4] in[5] in[6] in[7]
+ ctrl[0] ctrl[1] ctrl[2] out[0] out[1] out[2] out[3] out[4] out[5] out[6] out[7]
XNAND2X1_10 INVX1_11/A ctrl[0] gnd OAI21X1_11/C vdd NAND2X1
XNAND2X1_21 in[7] ctrl[2] gnd OAI21X1_22/C vdd NAND2X1
XOAI21X1_19 ctrl[2] INVX1_18/Y OAI21X1_19/C gnd INVX1_2/A vdd OAI21X1
XFILL_0_0_0 gnd vdd FILL
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XNAND2X1_22 gnd ctrl[2] gnd OAI21X1_23/C vdd NAND2X1
XNAND2X1_11 INVX1_12/A ctrl[0] gnd OAI21X1_12/C vdd NAND2X1
XFILL_0_0_1 gnd vdd FILL
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XNAND2X1_23 gnd ctrl[2] gnd OAI21X1_24/C vdd NAND2X1
XNAND2X1_12 INVX1_13/A ctrl[0] gnd NAND2X1_12/Y vdd NAND2X1
XFILL_0_0_2 gnd vdd FILL
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XNAND2X1_24 gnd ctrl[2] gnd OAI21X1_1/C vdd NAND2X1
XNAND2X1_13 INVX1_14/A ctrl[0] gnd NAND2X1_13/Y vdd NAND2X1
XFILL_3_0_0 gnd vdd FILL
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XNAND2X1_14 INVX1_15/A ctrl[0] gnd OAI21X1_15/C vdd NAND2X1
XFILL_3_0_1 gnd vdd FILL
XNAND2X1_15 INVX1_16/A ctrl[0] gnd OAI21X1_16/C vdd NAND2X1
XFILL_3_0_2 gnd vdd FILL
XNAND2X1_16 INVX1_17/A ctrl[0] gnd OAI21X1_17/C vdd NAND2X1
XFILL_1_1_0 gnd vdd FILL
XFILL_1_1_1 gnd vdd FILL
XNAND2X1_17 gnd ctrl[0] gnd NAND2X1_17/Y vdd NAND2X1
XNAND2X1_18 in[4] ctrl[2] gnd OAI21X1_19/C vdd NAND2X1
XFILL_1_1_2 gnd vdd FILL
XOAI21X1_1 ctrl[2] INVX1_24/Y OAI21X1_1/C gnd INVX1_8/A vdd OAI21X1
XNAND2X1_19 in[5] ctrl[2] gnd NAND2X1_19/Y vdd NAND2X1
XOAI21X1_2 ctrl[2] INVX1_1/Y NAND2X1_1/Y gnd INVX1_9/A vdd OAI21X1
XOAI21X1_3 ctrl[1] INVX1_2/Y OAI21X1_3/C gnd INVX1_10/A vdd OAI21X1
XBUFX2_1 BUFX2_1/A gnd out[0] vdd BUFX2
XOAI21X1_4 ctrl[1] INVX1_3/Y OAI21X1_4/C gnd INVX1_11/A vdd OAI21X1
XBUFX2_2 BUFX2_2/A gnd out[1] vdd BUFX2
XOAI21X1_5 ctrl[1] INVX1_4/Y NAND2X1_4/Y gnd INVX1_12/A vdd OAI21X1
XBUFX2_3 BUFX2_3/A gnd out[2] vdd BUFX2
XOAI21X1_6 ctrl[1] INVX1_5/Y OAI21X1_6/C gnd INVX1_13/A vdd OAI21X1
XFILL_2_0_0 gnd vdd FILL
XBUFX2_4 BUFX2_4/A gnd out[3] vdd BUFX2
XOAI21X1_7 ctrl[1] INVX1_6/Y NAND2X1_6/Y gnd INVX1_14/A vdd OAI21X1
XFILL_2_0_1 gnd vdd FILL
XBUFX2_5 BUFX2_5/A gnd out[4] vdd BUFX2
XOAI21X1_8 ctrl[1] INVX1_7/Y OAI21X1_8/C gnd INVX1_15/A vdd OAI21X1
XFILL_2_0_2 gnd vdd FILL
XFILL_0_1_0 gnd vdd FILL
XBUFX2_6 BUFX2_6/A gnd out[5] vdd BUFX2
XNAND2X1_1 gnd ctrl[2] gnd NAND2X1_1/Y vdd NAND2X1
XOAI21X1_9 ctrl[1] INVX1_8/Y OAI21X1_9/C gnd INVX1_16/A vdd OAI21X1
XNAND2X1_2 INVX1_4/A ctrl[1] gnd OAI21X1_3/C vdd NAND2X1
XFILL_0_1_1 gnd vdd FILL
XBUFX2_7 BUFX2_7/A gnd out[6] vdd BUFX2
XFILL_0_1_2 gnd vdd FILL
XBUFX2_8 BUFX2_8/A gnd out[7] vdd BUFX2
XNAND2X1_3 INVX1_5/A ctrl[1] gnd OAI21X1_4/C vdd NAND2X1
XFILL_3_1_0 gnd vdd FILL
XNAND2X1_4 INVX1_6/A ctrl[1] gnd NAND2X1_4/Y vdd NAND2X1
XFILL_3_1_1 gnd vdd FILL
XNAND2X1_5 INVX1_7/A ctrl[1] gnd OAI21X1_6/C vdd NAND2X1
XINVX1_20 in[2] gnd INVX1_20/Y vdd INVX1
XFILL_3_1_2 gnd vdd FILL
XINVX1_10 INVX1_10/A gnd INVX1_10/Y vdd INVX1
XNAND2X1_6 INVX1_8/A ctrl[1] gnd NAND2X1_6/Y vdd NAND2X1
XINVX1_21 in[3] gnd INVX1_21/Y vdd INVX1
XNAND2X1_7 INVX1_9/A ctrl[1] gnd OAI21X1_8/C vdd NAND2X1
XINVX1_22 in[4] gnd INVX1_22/Y vdd INVX1
XINVX1_11 INVX1_11/A gnd INVX1_11/Y vdd INVX1
XNAND2X1_8 gnd ctrl[1] gnd OAI21X1_9/C vdd NAND2X1
XINVX1_23 in[5] gnd INVX1_23/Y vdd INVX1
XINVX1_12 INVX1_12/A gnd INVX1_12/Y vdd INVX1
XINVX1_24 in[6] gnd INVX1_24/Y vdd INVX1
XINVX1_13 INVX1_13/A gnd INVX1_13/Y vdd INVX1
XNAND2X1_9 gnd ctrl[1] gnd NAND2X1_9/Y vdd NAND2X1
XFILL_1_0_0 gnd vdd FILL
XINVX1_14 INVX1_14/A gnd INVX1_14/Y vdd INVX1
XOAI21X1_20 ctrl[2] INVX1_19/Y NAND2X1_19/Y gnd INVX1_3/A vdd OAI21X1
XFILL_1_0_1 gnd vdd FILL
XINVX1_15 INVX1_15/A gnd INVX1_15/Y vdd INVX1
XOAI21X1_10 ctrl[1] INVX1_9/Y NAND2X1_9/Y gnd INVX1_17/A vdd OAI21X1
XOAI21X1_21 ctrl[2] INVX1_20/Y NAND2X1_20/Y gnd INVX1_4/A vdd OAI21X1
XFILL_1_0_2 gnd vdd FILL
XINVX1_16 INVX1_16/A gnd INVX1_16/Y vdd INVX1
XOAI21X1_11 ctrl[0] INVX1_10/Y OAI21X1_11/C gnd BUFX2_1/A vdd OAI21X1
XOAI21X1_22 ctrl[2] INVX1_21/Y OAI21X1_22/C gnd INVX1_5/A vdd OAI21X1
XINVX1_17 INVX1_17/A gnd INVX1_17/Y vdd INVX1
XOAI21X1_23 ctrl[2] INVX1_22/Y OAI21X1_23/C gnd INVX1_6/A vdd OAI21X1
XOAI21X1_12 ctrl[0] INVX1_11/Y OAI21X1_12/C gnd BUFX2_2/A vdd OAI21X1
XINVX1_18 in[0] gnd INVX1_18/Y vdd INVX1
XOAI21X1_24 ctrl[2] INVX1_23/Y OAI21X1_24/C gnd INVX1_7/A vdd OAI21X1
XOAI21X1_13 ctrl[0] INVX1_12/Y NAND2X1_12/Y gnd BUFX2_3/A vdd OAI21X1
XFILL_2_1_0 gnd vdd FILL
XINVX1_19 in[1] gnd INVX1_19/Y vdd INVX1
XOAI21X1_14 ctrl[0] INVX1_13/Y NAND2X1_13/Y gnd BUFX2_4/A vdd OAI21X1
XINVX1_1 in[7] gnd INVX1_1/Y vdd INVX1
XFILL_2_1_1 gnd vdd FILL
XOAI21X1_15 ctrl[0] INVX1_14/Y OAI21X1_15/C gnd BUFX2_5/A vdd OAI21X1
XINVX1_2 INVX1_2/A gnd INVX1_2/Y vdd INVX1
XFILL_2_1_2 gnd vdd FILL
XOAI21X1_16 ctrl[0] INVX1_15/Y OAI21X1_16/C gnd BUFX2_6/A vdd OAI21X1
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XOAI21X1_17 ctrl[0] INVX1_16/Y OAI21X1_17/C gnd BUFX2_7/A vdd OAI21X1
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XNAND2X1_20 in[6] ctrl[2] gnd NAND2X1_20/Y vdd NAND2X1
XOAI21X1_18 ctrl[0] INVX1_17/Y NAND2X1_17/Y gnd BUFX2_8/A vdd OAI21X1
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
.ends

