VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO barrel_shifter_8bit
  CLASS BLOCK ;
  FOREIGN barrel_shifter_8bit ;
  ORIGIN 1.900 4.000 ;
  SIZE 111.000 BY 88.300 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.400 80.400 106.800 81.600 ;
        RECT 1.200 75.800 2.000 80.400 ;
        RECT 4.400 71.800 5.200 80.400 ;
        RECT 8.600 75.800 9.400 80.400 ;
        RECT 10.800 75.800 11.600 80.400 ;
        RECT 14.000 71.800 14.800 80.400 ;
        RECT 18.200 75.800 19.000 80.400 ;
        RECT 20.400 75.800 21.200 80.400 ;
        RECT 23.600 75.800 24.400 80.400 ;
        RECT 31.600 73.000 32.400 80.400 ;
        RECT 36.400 75.800 37.200 80.400 ;
        RECT 38.000 71.800 38.800 80.400 ;
        RECT 42.200 75.800 43.000 80.400 ;
        RECT 44.400 75.800 45.200 80.400 ;
        RECT 47.600 75.800 48.400 80.400 ;
        RECT 49.200 75.800 50.000 80.400 ;
        RECT 52.400 71.800 53.200 80.400 ;
        RECT 56.600 75.800 57.400 80.400 ;
        RECT 58.800 75.800 59.600 80.400 ;
        RECT 62.000 71.800 62.800 80.400 ;
        RECT 66.200 75.800 67.000 80.400 ;
        RECT 70.000 73.000 70.800 80.400 ;
        RECT 78.000 75.800 78.800 80.400 ;
        RECT 81.200 75.800 82.000 80.400 ;
        RECT 82.800 75.800 83.600 80.400 ;
        RECT 86.000 71.800 86.800 80.400 ;
        RECT 90.200 75.800 91.000 80.400 ;
        RECT 92.400 75.800 93.200 80.400 ;
        RECT 95.600 75.800 96.400 80.400 ;
        RECT 97.200 75.800 98.000 80.400 ;
        RECT 101.000 75.800 101.800 80.400 ;
        RECT 105.200 71.800 106.000 80.400 ;
        RECT 1.200 41.600 2.000 46.200 ;
        RECT 4.400 41.600 5.200 46.200 ;
        RECT 6.000 41.600 6.800 46.200 ;
        RECT 9.200 41.600 10.000 46.200 ;
        RECT 12.400 41.600 13.200 46.200 ;
        RECT 14.000 41.600 14.800 46.200 ;
        RECT 17.200 41.600 18.000 50.200 ;
        RECT 21.400 41.600 22.200 46.200 ;
        RECT 23.600 41.600 24.400 46.200 ;
        RECT 26.800 41.600 27.600 46.200 ;
        RECT 33.200 41.600 34.000 50.200 ;
        RECT 37.400 41.600 38.200 46.200 ;
        RECT 39.600 41.600 40.400 46.200 ;
        RECT 42.800 41.600 43.600 46.200 ;
        RECT 44.400 41.600 45.200 46.200 ;
        RECT 47.600 41.600 48.400 46.200 ;
        RECT 50.800 41.600 51.600 46.200 ;
        RECT 52.400 41.600 53.200 50.200 ;
        RECT 56.600 41.600 57.400 46.200 ;
        RECT 58.800 41.600 59.600 46.200 ;
        RECT 62.000 41.600 62.800 46.200 ;
        RECT 63.600 41.600 64.400 46.200 ;
        RECT 66.800 41.600 67.600 46.200 ;
        RECT 68.400 41.600 69.200 46.200 ;
        RECT 71.600 41.600 72.400 46.200 ;
        RECT 80.200 41.600 81.000 46.200 ;
        RECT 84.400 41.600 85.200 50.200 ;
        RECT 86.000 41.600 86.800 46.200 ;
        RECT 89.200 41.600 90.000 46.200 ;
        RECT 90.800 41.600 91.600 46.200 ;
        RECT 94.000 41.600 94.800 46.200 ;
        RECT 96.200 41.600 97.000 46.200 ;
        RECT 100.400 41.600 101.200 50.200 ;
        RECT 103.600 41.600 104.400 49.000 ;
        RECT 0.400 40.400 106.800 41.600 ;
        RECT 1.200 35.800 2.000 40.400 ;
        RECT 6.000 33.000 6.800 40.400 ;
        RECT 9.800 35.800 10.600 40.400 ;
        RECT 14.000 31.800 14.800 40.400 ;
        RECT 17.200 35.800 18.000 40.400 ;
        RECT 18.800 35.800 19.600 40.400 ;
        RECT 22.000 35.800 22.800 40.400 ;
        RECT 28.400 31.800 29.200 40.400 ;
        RECT 32.600 35.800 33.400 40.400 ;
        RECT 34.800 35.800 35.600 40.400 ;
        RECT 38.000 31.800 38.800 40.400 ;
        RECT 42.200 35.800 43.000 40.400 ;
        RECT 44.400 35.800 45.200 40.400 ;
        RECT 47.600 35.800 48.400 40.400 ;
        RECT 49.200 35.800 50.000 40.400 ;
        RECT 52.400 35.800 53.200 40.400 ;
        RECT 54.000 35.800 54.800 40.400 ;
        RECT 57.200 31.800 58.000 40.400 ;
        RECT 61.400 35.800 62.200 40.400 ;
        RECT 63.600 35.800 64.400 40.400 ;
        RECT 66.800 35.800 67.600 40.400 ;
        RECT 68.400 35.800 69.200 40.400 ;
        RECT 71.600 35.800 72.400 40.400 ;
        RECT 78.000 35.800 78.800 40.400 ;
        RECT 81.200 31.800 82.000 40.400 ;
        RECT 85.400 35.800 86.200 40.400 ;
        RECT 87.600 35.800 88.400 40.400 ;
        RECT 90.800 35.800 91.600 40.400 ;
        RECT 92.400 35.800 93.200 40.400 ;
        RECT 95.600 35.800 96.400 40.400 ;
        RECT 98.800 33.000 99.600 40.400 ;
        RECT 103.600 33.000 104.400 40.400 ;
        RECT 1.200 1.600 2.000 6.200 ;
        RECT 4.400 1.600 5.200 10.200 ;
        RECT 8.600 1.600 9.400 6.200 ;
        RECT 10.800 1.600 11.600 6.200 ;
        RECT 14.000 1.600 14.800 10.200 ;
        RECT 18.200 1.600 19.000 6.200 ;
        RECT 20.400 1.600 21.200 6.200 ;
        RECT 23.600 1.600 24.400 6.200 ;
        RECT 30.000 1.600 30.800 6.200 ;
        RECT 33.200 1.600 34.000 6.200 ;
        RECT 36.400 1.600 37.200 6.200 ;
        RECT 38.000 1.600 38.800 10.200 ;
        RECT 42.200 1.600 43.000 6.200 ;
        RECT 44.400 1.600 45.200 6.200 ;
        RECT 47.600 1.600 48.400 6.200 ;
        RECT 49.200 1.600 50.000 6.200 ;
        RECT 52.400 1.600 53.200 10.200 ;
        RECT 56.600 1.600 57.400 6.200 ;
        RECT 58.800 1.600 59.600 6.200 ;
        RECT 62.000 1.600 62.800 6.200 ;
        RECT 63.600 1.600 64.400 6.200 ;
        RECT 67.400 1.600 68.200 6.200 ;
        RECT 71.600 1.600 72.400 10.200 ;
        RECT 78.600 1.600 79.400 6.200 ;
        RECT 82.800 1.600 83.600 10.200 ;
        RECT 86.000 1.600 86.800 6.200 ;
        RECT 89.200 1.600 90.000 9.000 ;
        RECT 92.400 1.600 93.200 6.200 ;
        RECT 96.200 1.600 97.000 6.200 ;
        RECT 100.400 1.600 101.200 10.200 ;
        RECT 103.600 1.600 104.400 9.000 ;
        RECT 0.400 0.400 106.800 1.600 ;
      LAYER via1 ;
        RECT 25.400 80.600 26.200 81.400 ;
        RECT 26.800 80.600 27.600 81.400 ;
        RECT 28.200 80.600 29.000 81.400 ;
        RECT 25.400 40.600 26.200 41.400 ;
        RECT 26.800 40.600 27.600 41.400 ;
        RECT 28.200 40.600 29.000 41.400 ;
        RECT 25.400 0.600 26.200 1.400 ;
        RECT 26.800 0.600 27.600 1.400 ;
        RECT 28.200 0.600 29.000 1.400 ;
      LAYER metal2 ;
        RECT 24.800 80.600 29.600 81.400 ;
        RECT 24.800 40.600 29.600 41.400 ;
        RECT 24.800 0.600 29.600 1.400 ;
      LAYER via2 ;
        RECT 25.400 80.600 26.200 81.400 ;
        RECT 26.800 80.600 27.600 81.400 ;
        RECT 28.200 80.600 29.000 81.400 ;
        RECT 25.400 40.600 26.200 41.400 ;
        RECT 26.800 40.600 27.600 41.400 ;
        RECT 28.200 40.600 29.000 41.400 ;
        RECT 25.400 0.600 26.200 1.400 ;
        RECT 26.800 0.600 27.600 1.400 ;
        RECT 28.200 0.600 29.000 1.400 ;
      LAYER metal3 ;
        RECT 24.800 80.400 29.600 81.600 ;
        RECT 24.800 40.400 29.600 41.600 ;
        RECT 24.800 0.400 29.600 1.600 ;
      LAYER via3 ;
        RECT 25.200 80.600 26.000 81.400 ;
        RECT 26.800 80.600 27.600 81.400 ;
        RECT 28.400 80.600 29.200 81.400 ;
        RECT 25.200 40.600 26.000 41.400 ;
        RECT 26.800 40.600 27.600 41.400 ;
        RECT 28.400 40.600 29.200 41.400 ;
        RECT 25.200 0.600 26.000 1.400 ;
        RECT 26.800 0.600 27.600 1.400 ;
        RECT 28.400 0.600 29.200 1.400 ;
      LAYER metal4 ;
        RECT 24.800 -4.000 29.600 84.000 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 1.200 61.600 2.000 64.200 ;
        RECT 6.000 61.600 6.800 65.400 ;
        RECT 10.800 61.600 11.600 64.200 ;
        RECT 15.600 61.600 16.400 65.400 ;
        RECT 23.600 61.600 24.400 66.200 ;
        RECT 31.600 61.600 32.400 66.200 ;
        RECT 36.400 61.600 37.200 64.200 ;
        RECT 39.600 61.600 40.400 65.400 ;
        RECT 47.600 61.600 48.400 66.200 ;
        RECT 49.200 61.600 50.000 64.200 ;
        RECT 54.000 61.600 54.800 65.400 ;
        RECT 58.800 61.600 59.600 64.200 ;
        RECT 63.600 61.600 64.400 65.400 ;
        RECT 70.000 61.600 70.800 66.200 ;
        RECT 78.000 61.600 78.800 66.200 ;
        RECT 82.800 61.600 83.600 64.200 ;
        RECT 87.600 61.600 88.400 65.400 ;
        RECT 95.600 61.600 96.400 66.200 ;
        RECT 97.200 61.600 98.000 64.200 ;
        RECT 103.600 61.600 104.400 65.400 ;
        RECT 0.400 60.400 106.800 61.600 ;
        RECT 1.200 55.800 2.000 60.400 ;
        RECT 6.000 57.800 6.800 60.400 ;
        RECT 12.400 55.800 13.200 60.400 ;
        RECT 14.000 57.800 14.800 60.400 ;
        RECT 18.800 56.600 19.600 60.400 ;
        RECT 26.800 55.800 27.600 60.400 ;
        RECT 34.800 56.600 35.600 60.400 ;
        RECT 42.800 55.800 43.600 60.400 ;
        RECT 44.400 57.800 45.200 60.400 ;
        RECT 47.600 55.800 48.400 60.400 ;
        RECT 54.000 56.600 54.800 60.400 ;
        RECT 62.000 55.800 62.800 60.400 ;
        RECT 63.600 55.800 64.400 60.400 ;
        RECT 68.400 57.800 69.200 60.400 ;
        RECT 71.600 57.800 72.400 60.400 ;
        RECT 82.800 56.600 83.600 60.400 ;
        RECT 89.200 55.800 90.000 60.400 ;
        RECT 90.800 55.800 91.600 60.400 ;
        RECT 98.800 56.600 99.600 60.400 ;
        RECT 103.600 55.800 104.400 60.400 ;
        RECT 47.700 55.200 48.300 55.800 ;
        RECT 42.800 53.600 43.600 55.200 ;
        RECT 47.600 53.600 48.400 55.200 ;
        RECT 89.200 53.600 90.000 55.200 ;
        RECT 90.800 53.600 91.600 55.200 ;
        RECT 47.600 26.800 48.400 28.400 ;
        RECT 49.200 26.800 50.000 28.400 ;
        RECT 66.800 26.800 67.600 28.400 ;
        RECT 1.200 21.600 2.000 24.200 ;
        RECT 6.000 21.600 6.800 26.200 ;
        RECT 12.400 21.600 13.200 25.400 ;
        RECT 17.200 21.600 18.000 24.200 ;
        RECT 22.000 21.600 22.800 26.200 ;
        RECT 30.000 21.600 30.800 25.400 ;
        RECT 34.800 21.600 35.600 24.200 ;
        RECT 39.600 21.600 40.400 25.400 ;
        RECT 47.600 21.600 48.400 26.200 ;
        RECT 49.200 21.600 50.000 26.200 ;
        RECT 54.000 21.600 54.800 24.200 ;
        RECT 58.800 21.600 59.600 25.400 ;
        RECT 66.800 21.600 67.600 26.200 ;
        RECT 68.400 21.600 69.200 26.200 ;
        RECT 78.000 21.600 78.800 24.200 ;
        RECT 82.800 21.600 83.600 25.400 ;
        RECT 87.600 21.600 88.400 26.200 ;
        RECT 92.400 21.600 93.200 26.200 ;
        RECT 98.800 21.600 99.600 26.200 ;
        RECT 103.600 21.600 104.400 26.200 ;
        RECT 0.400 20.400 106.800 21.600 ;
        RECT 1.200 17.800 2.000 20.400 ;
        RECT 6.000 16.600 6.800 20.400 ;
        RECT 10.800 17.800 11.600 20.400 ;
        RECT 15.600 16.600 16.400 20.400 ;
        RECT 23.600 15.800 24.400 20.400 ;
        RECT 30.000 17.800 30.800 20.400 ;
        RECT 36.400 15.800 37.200 20.400 ;
        RECT 39.600 16.600 40.400 20.400 ;
        RECT 47.600 15.800 48.400 20.400 ;
        RECT 49.200 17.800 50.000 20.400 ;
        RECT 54.000 16.600 54.800 20.400 ;
        RECT 58.800 15.800 59.600 20.400 ;
        RECT 63.600 17.800 64.400 20.400 ;
        RECT 70.000 16.600 70.800 20.400 ;
        RECT 81.200 16.600 82.000 20.400 ;
        RECT 86.000 17.800 86.800 20.400 ;
        RECT 89.200 15.800 90.000 20.400 ;
        RECT 92.400 17.800 93.200 20.400 ;
        RECT 98.800 16.600 99.600 20.400 ;
        RECT 103.600 15.800 104.400 20.400 ;
      LAYER via1 ;
        RECT 73.400 60.600 74.200 61.400 ;
        RECT 74.800 60.600 75.600 61.400 ;
        RECT 76.200 60.600 77.000 61.400 ;
        RECT 42.800 57.600 43.600 58.400 ;
        RECT 89.200 57.600 90.000 58.400 ;
        RECT 90.800 57.600 91.600 58.400 ;
        RECT 47.600 27.600 48.400 28.400 ;
        RECT 49.200 27.600 50.000 28.400 ;
        RECT 66.800 27.600 67.600 28.400 ;
        RECT 47.600 23.600 48.400 24.400 ;
        RECT 49.200 23.600 50.000 24.400 ;
        RECT 66.800 23.600 67.600 24.400 ;
        RECT 73.400 20.600 74.200 21.400 ;
        RECT 74.800 20.600 75.600 21.400 ;
        RECT 76.200 20.600 77.000 21.400 ;
      LAYER metal2 ;
        RECT 72.800 60.600 77.600 61.400 ;
        RECT 42.800 57.600 43.600 58.400 ;
        RECT 89.200 57.600 90.000 58.400 ;
        RECT 90.800 57.600 91.600 58.400 ;
        RECT 42.900 54.400 43.500 57.600 ;
        RECT 89.300 54.400 89.900 57.600 ;
        RECT 90.900 54.400 91.500 57.600 ;
        RECT 42.800 53.600 43.600 54.400 ;
        RECT 89.200 53.600 90.000 54.400 ;
        RECT 90.800 53.600 91.600 54.400 ;
        RECT 47.600 27.600 48.400 28.400 ;
        RECT 49.200 27.600 50.000 28.400 ;
        RECT 66.800 27.600 67.600 28.400 ;
        RECT 47.700 24.400 48.300 27.600 ;
        RECT 49.300 24.400 49.900 27.600 ;
        RECT 66.900 24.400 67.500 27.600 ;
        RECT 47.600 23.600 48.400 24.400 ;
        RECT 49.200 23.600 50.000 24.400 ;
        RECT 66.800 23.600 67.600 24.400 ;
        RECT 72.800 20.600 77.600 21.400 ;
      LAYER via2 ;
        RECT 73.400 60.600 74.200 61.400 ;
        RECT 74.800 60.600 75.600 61.400 ;
        RECT 76.200 60.600 77.000 61.400 ;
        RECT 73.400 20.600 74.200 21.400 ;
        RECT 74.800 20.600 75.600 21.400 ;
        RECT 76.200 20.600 77.000 21.400 ;
      LAYER metal3 ;
        RECT 72.800 60.400 77.600 61.600 ;
        RECT 72.800 20.400 77.600 21.600 ;
      LAYER via3 ;
        RECT 73.200 60.600 74.000 61.400 ;
        RECT 74.800 60.600 75.600 61.400 ;
        RECT 76.400 60.600 77.200 61.400 ;
        RECT 73.200 20.600 74.000 21.400 ;
        RECT 74.800 20.600 75.600 21.400 ;
        RECT 76.400 20.600 77.200 21.400 ;
      LAYER metal4 ;
        RECT 72.800 -4.000 77.600 84.000 ;
    END
  END gnd
  PIN in[0]
    PORT
      LAYER metal1 ;
        RECT 1.200 15.600 2.000 17.200 ;
      LAYER metal2 ;
        RECT 1.200 15.600 2.000 16.400 ;
        RECT 1.300 10.400 1.900 15.600 ;
        RECT 1.200 9.600 2.000 10.400 ;
      LAYER metal3 ;
        RECT 1.200 10.300 2.000 10.400 ;
        RECT -1.900 9.700 2.000 10.300 ;
        RECT 1.200 9.600 2.000 9.700 ;
    END
  END in[0]
  PIN in[1]
    PORT
      LAYER metal1 ;
        RECT 1.200 64.800 2.000 66.400 ;
      LAYER via1 ;
        RECT 1.200 65.600 2.000 66.400 ;
      LAYER metal2 ;
        RECT 1.200 69.600 2.000 70.400 ;
        RECT 1.300 66.400 1.900 69.600 ;
        RECT 1.200 65.600 2.000 66.400 ;
      LAYER metal3 ;
        RECT 1.200 70.300 2.000 70.400 ;
        RECT -1.900 69.700 2.000 70.300 ;
        RECT 1.200 69.600 2.000 69.700 ;
    END
  END in[1]
  PIN in[2]
    PORT
      LAYER metal1 ;
        RECT 1.200 24.800 2.000 26.400 ;
      LAYER via1 ;
        RECT 1.200 25.600 2.000 26.400 ;
      LAYER metal2 ;
        RECT 1.200 27.600 2.000 28.400 ;
        RECT 1.300 26.400 1.900 27.600 ;
        RECT 1.200 25.600 2.000 26.400 ;
      LAYER metal3 ;
        RECT 1.200 28.300 2.000 28.400 ;
        RECT -1.900 27.700 2.000 28.300 ;
        RECT 1.200 27.600 2.000 27.700 ;
    END
  END in[2]
  PIN in[3]
    PORT
      LAYER metal1 ;
        RECT 36.400 64.800 37.200 66.400 ;
      LAYER via1 ;
        RECT 36.400 65.600 37.200 66.400 ;
      LAYER metal2 ;
        RECT 34.900 83.700 37.100 84.300 ;
        RECT 36.500 66.400 37.100 83.700 ;
        RECT 36.400 65.600 37.200 66.400 ;
    END
  END in[3]
  PIN in[4]
    PORT
      LAYER metal1 ;
        RECT 30.000 15.600 30.800 17.200 ;
        RECT 23.600 14.300 24.400 15.200 ;
        RECT 30.100 14.400 30.700 15.600 ;
        RECT 30.000 14.300 30.800 14.400 ;
        RECT 23.600 13.700 30.800 14.300 ;
        RECT 23.600 13.600 24.400 13.700 ;
        RECT 30.000 13.600 30.800 13.700 ;
      LAYER metal2 ;
        RECT 30.000 13.600 30.800 14.400 ;
        RECT 30.100 4.300 30.700 13.600 ;
        RECT 30.100 3.700 32.300 4.300 ;
        RECT 31.700 -1.700 32.300 3.700 ;
        RECT 30.100 -2.300 32.300 -1.700 ;
    END
  END in[4]
  PIN in[5]
    PORT
      LAYER metal1 ;
        RECT 6.000 55.600 6.800 57.200 ;
        RECT 1.200 53.600 2.000 55.200 ;
      LAYER metal2 ;
        RECT 1.200 55.600 2.000 56.400 ;
        RECT 6.000 55.600 6.800 56.400 ;
        RECT 1.300 54.400 1.900 55.600 ;
        RECT 1.200 53.600 2.000 54.400 ;
      LAYER metal3 ;
        RECT 1.200 56.300 2.000 56.400 ;
        RECT 6.000 56.300 6.800 56.400 ;
        RECT -1.900 55.700 6.800 56.300 ;
        RECT 1.200 55.600 2.000 55.700 ;
        RECT 6.000 55.600 6.800 55.700 ;
    END
  END in[5]
  PIN in[6]
    PORT
      LAYER metal1 ;
        RECT 49.200 15.600 50.000 17.200 ;
        RECT 36.400 13.600 37.200 15.200 ;
      LAYER metal2 ;
        RECT 36.400 17.600 37.200 18.400 ;
        RECT 49.200 17.600 50.000 18.400 ;
        RECT 36.500 14.400 37.100 17.600 ;
        RECT 49.300 16.400 49.900 17.600 ;
        RECT 49.200 15.600 50.000 16.400 ;
        RECT 36.400 13.600 37.200 14.400 ;
        RECT 36.500 -1.700 37.100 13.600 ;
        RECT 34.900 -2.300 37.100 -1.700 ;
      LAYER metal3 ;
        RECT 36.400 18.300 37.200 18.400 ;
        RECT 49.200 18.300 50.000 18.400 ;
        RECT 36.400 17.700 50.000 18.300 ;
        RECT 36.400 17.600 37.200 17.700 ;
        RECT 49.200 17.600 50.000 17.700 ;
    END
  END in[6]
  PIN in[7]
    PORT
      LAYER metal1 ;
        RECT 47.600 68.300 48.400 68.400 ;
        RECT 47.600 67.700 49.900 68.300 ;
        RECT 47.600 66.800 48.400 67.700 ;
        RECT 49.300 66.400 49.900 67.700 ;
        RECT 49.200 64.800 50.000 66.400 ;
      LAYER via1 ;
        RECT 47.600 67.600 48.400 68.400 ;
      LAYER metal2 ;
        RECT 47.700 68.400 48.300 84.300 ;
        RECT 47.600 67.600 48.400 68.400 ;
    END
  END in[7]
  PIN ctrl[0]
    PORT
      LAYER metal1 ;
        RECT 92.400 71.600 93.200 73.200 ;
        RECT 62.000 68.200 62.800 68.400 ;
        RECT 105.200 68.200 106.000 68.400 ;
        RECT 62.000 67.600 63.600 68.200 ;
        RECT 62.800 67.200 63.600 67.600 ;
        RECT 104.400 67.600 106.000 68.200 ;
        RECT 104.400 67.200 105.200 67.600 ;
        RECT 18.000 54.400 18.800 54.800 ;
        RECT 17.200 53.800 18.800 54.400 ;
        RECT 99.600 54.400 100.400 54.800 ;
        RECT 99.600 53.800 101.200 54.400 ;
        RECT 17.200 53.600 18.000 53.800 ;
        RECT 100.400 53.600 101.200 53.800 ;
        RECT 9.200 48.800 10.000 50.400 ;
        RECT 23.600 48.800 24.400 50.400 ;
        RECT 66.800 48.800 67.600 50.400 ;
        RECT 94.000 48.800 94.800 50.400 ;
        RECT 71.600 31.600 72.400 33.200 ;
        RECT 90.800 31.600 91.600 33.200 ;
        RECT 95.600 31.600 96.400 33.200 ;
        RECT 14.000 28.200 14.800 28.400 ;
        RECT 13.200 27.600 14.800 28.200 ;
        RECT 81.200 28.200 82.000 28.400 ;
        RECT 81.200 27.600 82.800 28.200 ;
        RECT 13.200 27.200 14.000 27.600 ;
        RECT 82.000 27.200 82.800 27.600 ;
        RECT 82.000 14.400 82.800 14.800 ;
        RECT 99.600 14.400 100.400 14.800 ;
        RECT 82.000 13.800 83.600 14.400 ;
        RECT 99.600 13.800 101.200 14.400 ;
        RECT 82.800 13.600 83.600 13.800 ;
        RECT 100.400 13.600 101.200 13.800 ;
      LAYER via1 ;
        RECT 105.200 67.600 106.000 68.400 ;
        RECT 9.200 49.600 10.000 50.400 ;
        RECT 23.600 49.600 24.400 50.400 ;
        RECT 66.800 49.600 67.600 50.400 ;
        RECT 94.000 49.600 94.800 50.400 ;
        RECT 14.000 27.600 14.800 28.400 ;
      LAYER metal2 ;
        RECT 92.400 71.600 93.200 72.400 ;
        RECT 105.200 71.600 106.000 72.400 ;
        RECT 105.300 68.400 105.900 71.600 ;
        RECT 62.000 68.300 62.800 68.400 ;
        RECT 60.500 67.700 62.800 68.300 ;
        RECT 9.200 53.600 10.000 54.400 ;
        RECT 14.000 53.600 14.800 54.400 ;
        RECT 17.200 53.600 18.000 54.400 ;
        RECT 23.600 53.600 24.400 54.400 ;
        RECT 9.300 50.400 9.900 53.600 ;
        RECT 9.200 49.600 10.000 50.400 ;
        RECT 14.100 28.400 14.700 53.600 ;
        RECT 23.700 52.400 24.300 53.600 ;
        RECT 60.500 52.400 61.100 67.700 ;
        RECT 62.000 67.600 62.800 67.700 ;
        RECT 100.400 67.600 101.200 68.400 ;
        RECT 105.200 67.600 106.000 68.400 ;
        RECT 100.500 54.400 101.100 67.600 ;
        RECT 94.000 53.600 94.800 54.400 ;
        RECT 100.400 53.600 101.200 54.400 ;
        RECT 23.600 51.600 24.400 52.400 ;
        RECT 60.400 51.600 61.200 52.400 ;
        RECT 66.800 51.600 67.600 52.400 ;
        RECT 71.600 51.600 72.400 52.400 ;
        RECT 23.700 50.400 24.300 51.600 ;
        RECT 66.900 50.400 67.500 51.600 ;
        RECT 23.600 49.600 24.400 50.400 ;
        RECT 66.800 49.600 67.600 50.400 ;
        RECT 71.700 32.400 72.300 51.600 ;
        RECT 94.100 50.400 94.700 53.600 ;
        RECT 94.000 49.600 94.800 50.400 ;
        RECT 94.100 46.300 94.700 49.600 ;
        RECT 94.100 45.700 96.300 46.300 ;
        RECT 95.700 32.400 96.300 45.700 ;
        RECT 71.600 31.600 72.400 32.400 ;
        RECT 90.800 31.600 91.600 32.400 ;
        RECT 95.600 31.600 96.400 32.400 ;
        RECT 71.700 30.400 72.300 31.600 ;
        RECT 90.900 30.400 91.500 31.600 ;
        RECT 95.700 30.400 96.300 31.600 ;
        RECT 71.600 29.600 72.400 30.400 ;
        RECT 81.200 29.600 82.000 30.400 ;
        RECT 82.800 29.600 83.600 30.400 ;
        RECT 90.800 29.600 91.600 30.400 ;
        RECT 95.600 29.600 96.400 30.400 ;
        RECT 81.300 28.400 81.900 29.600 ;
        RECT 14.000 27.600 14.800 28.400 ;
        RECT 81.200 27.600 82.000 28.400 ;
        RECT 82.900 14.400 83.500 29.600 ;
        RECT 95.700 14.400 96.300 29.600 ;
        RECT 82.800 13.600 83.600 14.400 ;
        RECT 95.600 13.600 96.400 14.400 ;
        RECT 100.400 13.600 101.200 14.400 ;
      LAYER metal3 ;
        RECT 92.400 72.300 93.200 72.400 ;
        RECT 105.200 72.300 106.000 72.400 ;
        RECT 92.400 71.700 106.000 72.300 ;
        RECT 92.400 71.600 93.200 71.700 ;
        RECT 105.200 71.600 106.000 71.700 ;
        RECT 100.400 68.300 101.200 68.400 ;
        RECT 105.200 68.300 106.000 68.400 ;
        RECT 100.400 67.700 109.100 68.300 ;
        RECT 100.400 67.600 101.200 67.700 ;
        RECT 105.200 67.600 106.000 67.700 ;
        RECT 9.200 54.300 10.000 54.400 ;
        RECT 14.000 54.300 14.800 54.400 ;
        RECT 17.200 54.300 18.000 54.400 ;
        RECT 23.600 54.300 24.400 54.400 ;
        RECT 9.200 53.700 24.400 54.300 ;
        RECT 9.200 53.600 10.000 53.700 ;
        RECT 14.000 53.600 14.800 53.700 ;
        RECT 17.200 53.600 18.000 53.700 ;
        RECT 23.600 53.600 24.400 53.700 ;
        RECT 94.000 54.300 94.800 54.400 ;
        RECT 100.400 54.300 101.200 54.400 ;
        RECT 94.000 53.700 101.200 54.300 ;
        RECT 94.000 53.600 94.800 53.700 ;
        RECT 100.400 53.600 101.200 53.700 ;
        RECT 23.600 52.300 24.400 52.400 ;
        RECT 60.400 52.300 61.200 52.400 ;
        RECT 66.800 52.300 67.600 52.400 ;
        RECT 71.600 52.300 72.400 52.400 ;
        RECT 23.600 51.700 72.400 52.300 ;
        RECT 23.600 51.600 24.400 51.700 ;
        RECT 60.400 51.600 61.200 51.700 ;
        RECT 66.800 51.600 67.600 51.700 ;
        RECT 71.600 51.600 72.400 51.700 ;
        RECT 71.600 30.300 72.400 30.400 ;
        RECT 81.200 30.300 82.000 30.400 ;
        RECT 82.800 30.300 83.600 30.400 ;
        RECT 90.800 30.300 91.600 30.400 ;
        RECT 95.600 30.300 96.400 30.400 ;
        RECT 71.600 29.700 96.400 30.300 ;
        RECT 71.600 29.600 72.400 29.700 ;
        RECT 81.200 29.600 82.000 29.700 ;
        RECT 82.800 29.600 83.600 29.700 ;
        RECT 90.800 29.600 91.600 29.700 ;
        RECT 95.600 29.600 96.400 29.700 ;
        RECT 95.600 14.300 96.400 14.400 ;
        RECT 100.400 14.300 101.200 14.400 ;
        RECT 95.600 13.700 101.200 14.300 ;
        RECT 95.600 13.600 96.400 13.700 ;
        RECT 100.400 13.600 101.200 13.700 ;
    END
  END ctrl[0]
  PIN ctrl[1]
    PORT
      LAYER metal1 ;
        RECT 20.400 71.600 21.200 73.200 ;
        RECT 81.200 71.600 82.000 73.200 ;
        RECT 14.000 68.200 14.800 68.400 ;
        RECT 86.000 68.200 86.800 68.400 ;
        RECT 14.000 67.600 15.600 68.200 ;
        RECT 86.000 67.600 87.600 68.200 ;
        RECT 14.800 67.200 15.600 67.600 ;
        RECT 86.800 67.200 87.600 67.600 ;
        RECT 53.200 54.400 54.000 54.800 ;
        RECT 52.400 53.800 54.000 54.400 ;
        RECT 83.600 54.400 84.400 54.800 ;
        RECT 83.600 54.300 85.200 54.400 ;
        RECT 86.000 54.300 86.800 54.400 ;
        RECT 83.600 53.800 86.800 54.300 ;
        RECT 52.400 53.600 53.200 53.800 ;
        RECT 84.400 53.700 86.800 53.800 ;
        RECT 84.400 53.600 85.200 53.700 ;
        RECT 86.000 53.600 86.800 53.700 ;
        RECT 58.800 48.800 59.600 50.400 ;
        RECT 86.000 48.800 86.800 50.400 ;
        RECT 18.800 31.600 19.600 33.200 ;
        RECT 63.600 31.600 64.400 33.200 ;
        RECT 38.000 28.200 38.800 28.400 ;
        RECT 57.200 28.200 58.000 28.400 ;
        RECT 38.000 27.600 39.600 28.200 ;
        RECT 57.200 27.600 58.800 28.200 ;
        RECT 38.800 27.200 39.600 27.600 ;
        RECT 58.000 27.200 58.800 27.600 ;
        RECT 14.800 14.400 15.600 14.800 ;
        RECT 14.000 13.800 15.600 14.400 ;
        RECT 70.800 14.400 71.600 14.800 ;
        RECT 70.800 13.800 72.400 14.400 ;
        RECT 14.000 13.600 14.800 13.800 ;
        RECT 71.600 13.600 72.400 13.800 ;
        RECT 44.400 8.800 45.200 10.400 ;
        RECT 62.000 8.800 62.800 10.400 ;
      LAYER via1 ;
        RECT 58.800 49.600 59.600 50.400 ;
        RECT 86.000 49.600 86.800 50.400 ;
        RECT 44.400 9.600 45.200 10.400 ;
        RECT 62.000 9.600 62.800 10.400 ;
      LAYER metal2 ;
        RECT 78.100 80.400 78.700 84.300 ;
        RECT 78.000 79.600 78.800 80.400 ;
        RECT 81.200 79.600 82.000 80.400 ;
        RECT 81.300 72.400 81.900 79.600 ;
        RECT 20.400 71.600 21.200 72.400 ;
        RECT 81.200 71.600 82.000 72.400 ;
        RECT 20.500 68.400 21.100 71.600 ;
        RECT 81.300 68.400 81.900 71.600 ;
        RECT 14.000 67.600 14.800 68.400 ;
        RECT 20.400 67.600 21.200 68.400 ;
        RECT 81.200 67.600 82.000 68.400 ;
        RECT 86.000 67.600 86.800 68.400 ;
        RECT 18.800 31.600 19.600 32.400 ;
        RECT 18.900 26.400 19.500 31.600 ;
        RECT 20.500 26.400 21.100 67.600 ;
        RECT 86.100 54.400 86.700 67.600 ;
        RECT 52.400 53.600 53.200 54.400 ;
        RECT 86.000 53.600 86.800 54.400 ;
        RECT 52.500 48.400 53.100 53.600 ;
        RECT 86.100 50.400 86.700 53.600 ;
        RECT 58.800 49.600 59.600 50.400 ;
        RECT 86.000 49.600 86.800 50.400 ;
        RECT 58.900 48.400 59.500 49.600 ;
        RECT 86.100 48.400 86.700 49.600 ;
        RECT 52.400 47.600 53.200 48.400 ;
        RECT 58.800 47.600 59.600 48.400 ;
        RECT 86.000 47.600 86.800 48.400 ;
        RECT 58.900 32.400 59.500 47.600 ;
        RECT 57.200 31.600 58.000 32.400 ;
        RECT 58.800 31.600 59.600 32.400 ;
        RECT 63.600 31.600 64.400 32.400 ;
        RECT 57.300 28.400 57.900 31.600 ;
        RECT 38.000 27.600 38.800 28.400 ;
        RECT 57.200 27.600 58.000 28.400 ;
        RECT 38.100 26.400 38.700 27.600 ;
        RECT 57.300 26.400 57.900 27.600 ;
        RECT 14.000 25.600 14.800 26.400 ;
        RECT 18.800 25.600 19.600 26.400 ;
        RECT 20.400 25.600 21.200 26.400 ;
        RECT 38.000 25.600 38.800 26.400 ;
        RECT 57.200 25.600 58.000 26.400 ;
        RECT 62.000 25.600 62.800 26.400 ;
        RECT 14.100 14.400 14.700 25.600 ;
        RECT 14.000 13.600 14.800 14.400 ;
        RECT 62.100 12.400 62.700 25.600 ;
        RECT 71.600 13.600 72.400 14.400 ;
        RECT 71.700 12.400 72.300 13.600 ;
        RECT 44.400 11.600 45.200 12.400 ;
        RECT 62.000 11.600 62.800 12.400 ;
        RECT 71.600 11.600 72.400 12.400 ;
        RECT 44.500 10.400 45.100 11.600 ;
        RECT 62.100 10.400 62.700 11.600 ;
        RECT 44.400 9.600 45.200 10.400 ;
        RECT 62.000 9.600 62.800 10.400 ;
      LAYER metal3 ;
        RECT 78.000 80.300 78.800 80.400 ;
        RECT 81.200 80.300 82.000 80.400 ;
        RECT 78.000 79.700 82.000 80.300 ;
        RECT 78.000 79.600 78.800 79.700 ;
        RECT 81.200 79.600 82.000 79.700 ;
        RECT 14.000 68.300 14.800 68.400 ;
        RECT 20.400 68.300 21.200 68.400 ;
        RECT 14.000 67.700 21.200 68.300 ;
        RECT 14.000 67.600 14.800 67.700 ;
        RECT 20.400 67.600 21.200 67.700 ;
        RECT 81.200 68.300 82.000 68.400 ;
        RECT 86.000 68.300 86.800 68.400 ;
        RECT 81.200 67.700 86.800 68.300 ;
        RECT 81.200 67.600 82.000 67.700 ;
        RECT 86.000 67.600 86.800 67.700 ;
        RECT 52.400 48.300 53.200 48.400 ;
        RECT 58.800 48.300 59.600 48.400 ;
        RECT 86.000 48.300 86.800 48.400 ;
        RECT 52.400 47.700 86.800 48.300 ;
        RECT 52.400 47.600 53.200 47.700 ;
        RECT 58.800 47.600 59.600 47.700 ;
        RECT 86.000 47.600 86.800 47.700 ;
        RECT 57.200 32.300 58.000 32.400 ;
        RECT 58.800 32.300 59.600 32.400 ;
        RECT 63.600 32.300 64.400 32.400 ;
        RECT 57.200 31.700 64.400 32.300 ;
        RECT 57.200 31.600 58.000 31.700 ;
        RECT 58.800 31.600 59.600 31.700 ;
        RECT 63.600 31.600 64.400 31.700 ;
        RECT 14.000 26.300 14.800 26.400 ;
        RECT 18.800 26.300 19.600 26.400 ;
        RECT 20.400 26.300 21.200 26.400 ;
        RECT 38.000 26.300 38.800 26.400 ;
        RECT 57.200 26.300 58.000 26.400 ;
        RECT 62.000 26.300 62.800 26.400 ;
        RECT 14.000 25.700 62.800 26.300 ;
        RECT 14.000 25.600 14.800 25.700 ;
        RECT 18.800 25.600 19.600 25.700 ;
        RECT 20.400 25.600 21.200 25.700 ;
        RECT 38.000 25.600 38.800 25.700 ;
        RECT 57.200 25.600 58.000 25.700 ;
        RECT 62.000 25.600 62.800 25.700 ;
        RECT 44.400 12.300 45.200 12.400 ;
        RECT 62.000 12.300 62.800 12.400 ;
        RECT 71.600 12.300 72.400 12.400 ;
        RECT 44.400 11.700 72.400 12.300 ;
        RECT 44.400 11.600 45.200 11.700 ;
        RECT 62.000 11.600 62.800 11.700 ;
        RECT 71.600 11.600 72.400 11.700 ;
    END
  END ctrl[1]
  PIN ctrl[2]
    PORT
      LAYER metal1 ;
        RECT 44.400 71.600 45.200 73.200 ;
        RECT 4.400 68.200 5.200 68.400 ;
        RECT 38.000 68.200 38.800 68.400 ;
        RECT 52.400 68.200 53.200 68.400 ;
        RECT 4.400 67.600 6.000 68.200 ;
        RECT 38.000 67.600 39.600 68.200 ;
        RECT 52.400 67.600 54.000 68.200 ;
        RECT 5.200 67.200 6.000 67.600 ;
        RECT 38.800 67.200 39.600 67.600 ;
        RECT 53.200 67.200 54.000 67.600 ;
        RECT 34.000 54.400 34.800 54.800 ;
        RECT 31.600 54.300 32.400 54.400 ;
        RECT 33.200 54.300 34.800 54.400 ;
        RECT 31.600 53.800 34.800 54.300 ;
        RECT 31.600 53.700 34.000 53.800 ;
        RECT 31.600 53.600 32.400 53.700 ;
        RECT 33.200 53.600 34.000 53.700 ;
        RECT 4.400 50.300 5.200 50.400 ;
        RECT 6.000 50.300 6.800 50.400 ;
        RECT 4.400 49.700 6.800 50.300 ;
        RECT 4.400 48.800 5.200 49.700 ;
        RECT 6.000 49.600 6.800 49.700 ;
        RECT 39.600 48.800 40.400 50.400 ;
        RECT 50.800 48.800 51.600 50.400 ;
        RECT 44.400 31.600 45.200 33.200 ;
        RECT 52.400 31.600 53.200 33.200 ;
        RECT 28.400 28.200 29.200 28.400 ;
        RECT 28.400 27.600 30.000 28.200 ;
        RECT 29.200 27.200 30.000 27.600 ;
        RECT 5.200 14.400 6.000 14.800 ;
        RECT 38.800 14.400 39.600 14.800 ;
        RECT 53.200 14.400 54.000 14.800 ;
        RECT 4.400 13.800 6.000 14.400 ;
        RECT 38.000 13.800 39.600 14.400 ;
        RECT 52.400 13.800 54.000 14.400 ;
        RECT 4.400 13.600 5.200 13.800 ;
        RECT 38.000 13.600 38.800 13.800 ;
        RECT 52.400 13.600 53.200 13.800 ;
        RECT 20.400 8.800 21.200 10.400 ;
        RECT 33.200 8.800 34.000 10.400 ;
      LAYER via1 ;
        RECT 39.600 49.600 40.400 50.400 ;
        RECT 50.800 49.600 51.600 50.400 ;
        RECT 20.400 9.600 21.200 10.400 ;
        RECT 33.200 9.600 34.000 10.400 ;
      LAYER metal2 ;
        RECT 39.600 71.600 40.400 72.400 ;
        RECT 44.400 71.600 45.200 72.400 ;
        RECT 4.400 67.600 5.200 68.400 ;
        RECT 38.000 68.300 38.800 68.400 ;
        RECT 39.700 68.300 40.300 71.600 ;
        RECT 44.500 68.400 45.100 71.600 ;
        RECT 38.000 67.700 40.300 68.300 ;
        RECT 38.000 67.600 38.800 67.700 ;
        RECT 4.500 52.400 5.100 67.600 ;
        RECT 31.600 53.600 32.400 54.400 ;
        RECT 4.400 51.600 5.200 52.400 ;
        RECT 6.000 51.600 6.800 52.400 ;
        RECT 6.100 50.400 6.700 51.600 ;
        RECT 31.700 50.400 32.300 53.600 ;
        RECT 39.700 50.400 40.300 67.700 ;
        RECT 44.400 67.600 45.200 68.400 ;
        RECT 52.400 67.600 53.200 68.400 ;
        RECT 6.000 49.600 6.800 50.400 ;
        RECT 31.600 49.600 32.400 50.400 ;
        RECT 39.600 49.600 40.400 50.400 ;
        RECT 50.800 49.600 51.600 50.400 ;
        RECT 6.100 14.400 6.700 49.600 ;
        RECT 31.700 32.400 32.300 49.600 ;
        RECT 50.900 32.400 51.500 49.600 ;
        RECT 28.400 31.600 29.200 32.400 ;
        RECT 31.600 31.600 32.400 32.400 ;
        RECT 44.400 31.600 45.200 32.400 ;
        RECT 50.800 31.600 51.600 32.400 ;
        RECT 52.400 31.600 53.200 32.400 ;
        RECT 28.500 28.400 29.100 31.600 ;
        RECT 28.400 27.600 29.200 28.400 ;
        RECT 52.500 14.400 53.100 31.600 ;
        RECT 4.400 13.600 5.200 14.400 ;
        RECT 6.000 13.600 6.800 14.400 ;
        RECT 20.400 13.600 21.200 14.400 ;
        RECT 33.200 13.600 34.000 14.400 ;
        RECT 38.000 13.600 38.800 14.400 ;
        RECT 52.400 13.600 53.200 14.400 ;
        RECT 20.500 10.400 21.100 13.600 ;
        RECT 33.300 10.400 33.900 13.600 ;
        RECT 20.400 9.600 21.200 10.400 ;
        RECT 33.200 9.600 34.000 10.400 ;
      LAYER metal3 ;
        RECT 39.600 72.300 40.400 72.400 ;
        RECT 44.400 72.300 45.200 72.400 ;
        RECT 39.600 71.700 45.200 72.300 ;
        RECT 39.600 71.600 40.400 71.700 ;
        RECT 44.400 71.600 45.200 71.700 ;
        RECT 44.400 68.300 45.200 68.400 ;
        RECT 52.400 68.300 53.200 68.400 ;
        RECT 44.400 67.700 53.200 68.300 ;
        RECT 44.400 67.600 45.200 67.700 ;
        RECT 52.400 67.600 53.200 67.700 ;
        RECT 4.400 52.300 5.200 52.400 ;
        RECT 6.000 52.300 6.800 52.400 ;
        RECT -1.900 51.700 6.800 52.300 ;
        RECT 4.400 51.600 5.200 51.700 ;
        RECT 6.000 51.600 6.800 51.700 ;
        RECT 31.600 50.300 32.400 50.400 ;
        RECT 39.600 50.300 40.400 50.400 ;
        RECT 31.600 49.700 40.400 50.300 ;
        RECT 31.600 49.600 32.400 49.700 ;
        RECT 39.600 49.600 40.400 49.700 ;
        RECT 28.400 32.300 29.200 32.400 ;
        RECT 31.600 32.300 32.400 32.400 ;
        RECT 44.400 32.300 45.200 32.400 ;
        RECT 50.800 32.300 51.600 32.400 ;
        RECT 52.400 32.300 53.200 32.400 ;
        RECT 28.400 31.700 53.200 32.300 ;
        RECT 28.400 31.600 29.200 31.700 ;
        RECT 31.600 31.600 32.400 31.700 ;
        RECT 44.400 31.600 45.200 31.700 ;
        RECT 50.800 31.600 51.600 31.700 ;
        RECT 52.400 31.600 53.200 31.700 ;
        RECT 4.400 14.300 5.200 14.400 ;
        RECT 6.000 14.300 6.800 14.400 ;
        RECT 20.400 14.300 21.200 14.400 ;
        RECT 33.200 14.300 34.000 14.400 ;
        RECT 38.000 14.300 38.800 14.400 ;
        RECT 52.400 14.300 53.200 14.400 ;
        RECT 4.400 13.700 53.200 14.300 ;
        RECT 4.400 13.600 5.200 13.700 ;
        RECT 6.000 13.600 6.800 13.700 ;
        RECT 20.400 13.600 21.200 13.700 ;
        RECT 33.200 13.600 34.000 13.700 ;
        RECT 38.000 13.600 38.800 13.700 ;
        RECT 52.400 13.600 53.200 13.700 ;
    END
  END ctrl[2]
  PIN out[0]
    PORT
      LAYER metal1 ;
        RECT 4.400 31.800 5.200 39.800 ;
        RECT 4.400 29.600 5.000 31.800 ;
        RECT 4.400 22.200 5.200 29.600 ;
      LAYER via1 ;
        RECT 4.400 33.600 5.200 34.400 ;
      LAYER metal2 ;
        RECT 4.400 33.600 5.200 34.400 ;
        RECT 4.500 32.400 5.100 33.600 ;
        RECT 4.400 31.600 5.200 32.400 ;
      LAYER metal3 ;
        RECT 4.400 32.300 5.200 32.400 ;
        RECT -1.900 31.700 5.200 32.300 ;
        RECT 4.400 31.600 5.200 31.700 ;
    END
  END out[0]
  PIN out[1]
    PORT
      LAYER metal1 ;
        RECT 33.200 71.800 34.000 79.800 ;
        RECT 33.400 69.600 34.000 71.800 ;
        RECT 33.200 62.200 34.000 69.600 ;
      LAYER via1 ;
        RECT 33.200 77.600 34.000 78.400 ;
      LAYER metal2 ;
        RECT 30.100 83.700 33.900 84.300 ;
        RECT 33.300 78.400 33.900 83.700 ;
        RECT 33.200 77.600 34.000 78.400 ;
    END
  END out[1]
  PIN out[2]
    PORT
      LAYER metal1 ;
        RECT 71.600 71.800 72.400 79.800 ;
        RECT 71.800 69.600 72.400 71.800 ;
        RECT 71.600 62.200 72.400 69.600 ;
      LAYER via1 ;
        RECT 71.600 77.600 72.400 78.400 ;
      LAYER metal2 ;
        RECT 70.100 83.700 72.300 84.300 ;
        RECT 71.700 78.400 72.300 83.700 ;
        RECT 71.600 77.600 72.400 78.400 ;
    END
  END out[2]
  PIN out[3]
    PORT
      LAYER metal1 ;
        RECT 105.200 52.400 106.000 59.800 ;
        RECT 105.400 50.200 106.000 52.400 ;
        RECT 105.200 42.200 106.000 50.200 ;
      LAYER via1 ;
        RECT 105.200 47.600 106.000 48.400 ;
      LAYER metal2 ;
        RECT 105.200 49.600 106.000 50.400 ;
        RECT 105.300 48.400 105.900 49.600 ;
        RECT 105.200 47.600 106.000 48.400 ;
      LAYER metal3 ;
        RECT 105.200 50.300 106.000 50.400 ;
        RECT 105.200 49.700 109.100 50.300 ;
        RECT 105.200 49.600 106.000 49.700 ;
    END
  END out[3]
  PIN out[4]
    PORT
      LAYER metal1 ;
        RECT 105.200 12.400 106.000 19.800 ;
        RECT 105.400 10.200 106.000 12.400 ;
        RECT 105.200 2.200 106.000 10.200 ;
      LAYER via1 ;
        RECT 105.200 7.600 106.000 8.400 ;
      LAYER metal2 ;
        RECT 105.200 9.600 106.000 10.400 ;
        RECT 105.300 8.400 105.900 9.600 ;
        RECT 105.200 7.600 106.000 8.400 ;
      LAYER metal3 ;
        RECT 105.200 10.300 106.000 10.400 ;
        RECT 105.200 9.700 109.100 10.300 ;
        RECT 105.200 9.600 106.000 9.700 ;
    END
  END out[4]
  PIN out[5]
    PORT
      LAYER metal1 ;
        RECT 90.800 12.400 91.600 19.800 ;
        RECT 91.000 10.200 91.600 12.400 ;
        RECT 90.800 2.200 91.600 10.200 ;
      LAYER via1 ;
        RECT 90.800 3.600 91.600 4.400 ;
      LAYER metal2 ;
        RECT 90.800 3.600 91.600 4.400 ;
        RECT 90.900 -1.700 91.500 3.600 ;
        RECT 89.300 -2.300 91.500 -1.700 ;
    END
  END out[5]
  PIN out[6]
    PORT
      LAYER metal1 ;
        RECT 100.400 31.800 101.200 39.800 ;
        RECT 100.600 29.600 101.200 31.800 ;
        RECT 100.400 22.200 101.200 29.600 ;
      LAYER via1 ;
        RECT 100.400 27.600 101.200 28.400 ;
      LAYER metal2 ;
        RECT 100.400 29.600 101.200 30.400 ;
        RECT 100.500 28.400 101.100 29.600 ;
        RECT 100.400 27.600 101.200 28.400 ;
      LAYER metal3 ;
        RECT 100.400 30.300 101.200 30.400 ;
        RECT 100.400 29.700 109.100 30.300 ;
        RECT 100.400 29.600 101.200 29.700 ;
    END
  END out[6]
  PIN out[7]
    PORT
      LAYER metal1 ;
        RECT 105.200 31.800 106.000 39.800 ;
        RECT 105.400 29.600 106.000 31.800 ;
        RECT 105.200 22.200 106.000 29.600 ;
      LAYER via1 ;
        RECT 105.200 33.600 106.000 34.400 ;
      LAYER metal2 ;
        RECT 105.200 33.600 106.000 34.400 ;
      LAYER metal3 ;
        RECT 105.200 34.300 106.000 34.400 ;
        RECT 105.200 33.700 109.100 34.300 ;
        RECT 105.200 33.600 106.000 33.700 ;
    END
  END out[7]
  OBS
      LAYER metal1 ;
        RECT 2.800 70.300 3.600 79.800 ;
        RECT 7.000 72.400 7.800 79.800 ;
        RECT 8.400 73.600 9.200 74.400 ;
        RECT 8.600 72.400 9.200 73.600 ;
        RECT 7.000 71.800 8.000 72.400 ;
        RECT 8.600 71.800 10.000 72.400 ;
        RECT 6.000 70.300 6.800 70.400 ;
        RECT 2.800 69.700 6.800 70.300 ;
        RECT 2.800 62.200 3.600 69.700 ;
        RECT 6.000 68.800 6.800 69.700 ;
        RECT 7.400 68.400 8.000 71.800 ;
        RECT 9.200 71.600 10.000 71.800 ;
        RECT 12.400 70.300 13.200 79.800 ;
        RECT 16.600 72.400 17.400 79.800 ;
        RECT 18.000 73.600 18.800 74.400 ;
        RECT 18.200 72.400 18.800 73.600 ;
        RECT 15.600 71.600 17.600 72.400 ;
        RECT 18.200 71.800 19.600 72.400 ;
        RECT 18.800 71.600 19.600 71.800 ;
        RECT 15.600 70.300 16.400 70.400 ;
        RECT 12.400 69.700 16.400 70.300 ;
        RECT 7.400 67.600 10.000 68.400 ;
        RECT 4.600 66.200 8.200 66.600 ;
        RECT 9.200 66.300 9.800 67.600 ;
        RECT 10.800 66.300 11.600 66.400 ;
        RECT 4.400 66.000 8.400 66.200 ;
        RECT 4.400 62.200 5.200 66.000 ;
        RECT 7.600 62.200 8.400 66.000 ;
        RECT 9.200 65.700 11.600 66.300 ;
        RECT 9.200 62.200 10.000 65.700 ;
        RECT 10.800 64.800 11.600 65.700 ;
        RECT 12.400 62.200 13.200 69.700 ;
        RECT 15.600 68.800 16.400 69.700 ;
        RECT 17.000 68.400 17.600 71.600 ;
        RECT 18.900 70.300 19.500 71.600 ;
        RECT 22.000 70.300 22.800 79.800 ;
        RECT 30.000 72.400 30.800 79.800 ;
        RECT 30.000 71.800 32.200 72.400 ;
        RECT 31.600 71.200 32.200 71.800 ;
        RECT 31.600 70.400 32.800 71.200 ;
        RECT 18.900 69.700 22.800 70.300 ;
        RECT 17.000 67.600 19.600 68.400 ;
        RECT 14.200 66.200 17.800 66.600 ;
        RECT 18.800 66.200 19.400 67.600 ;
        RECT 22.000 66.200 22.800 69.700 ;
        RECT 23.600 70.300 24.400 70.400 ;
        RECT 30.000 70.300 30.800 70.400 ;
        RECT 23.600 69.700 30.800 70.300 ;
        RECT 23.600 69.600 24.400 69.700 ;
        RECT 30.000 68.800 30.800 69.700 ;
        RECT 23.600 68.300 24.400 68.400 ;
        RECT 28.400 68.300 29.200 68.400 ;
        RECT 23.600 67.700 29.200 68.300 ;
        RECT 23.600 66.800 24.400 67.700 ;
        RECT 28.400 67.600 29.200 67.700 ;
        RECT 31.600 67.400 32.200 70.400 ;
        RECT 30.000 66.800 32.200 67.400 ;
        RECT 34.800 70.300 35.600 79.800 ;
        RECT 40.600 72.400 41.400 79.800 ;
        RECT 42.000 73.600 42.800 74.400 ;
        RECT 42.200 72.400 42.800 73.600 ;
        RECT 40.600 71.800 41.600 72.400 ;
        RECT 42.200 71.800 43.600 72.400 ;
        RECT 39.600 70.300 40.400 70.400 ;
        RECT 34.800 69.700 40.400 70.300 ;
        RECT 14.000 66.000 18.000 66.200 ;
        RECT 14.000 62.200 14.800 66.000 ;
        RECT 17.200 62.200 18.000 66.000 ;
        RECT 18.800 62.200 19.600 66.200 ;
        RECT 21.000 65.600 22.800 66.200 ;
        RECT 21.000 62.200 21.800 65.600 ;
        RECT 30.000 62.200 30.800 66.800 ;
        RECT 34.800 62.200 35.600 69.700 ;
        RECT 39.600 68.800 40.400 69.700 ;
        RECT 41.000 68.400 41.600 71.800 ;
        RECT 42.800 71.600 43.600 71.800 ;
        RECT 42.900 70.300 43.500 71.600 ;
        RECT 46.000 70.300 46.800 79.800 ;
        RECT 42.900 69.700 46.800 70.300 ;
        RECT 41.000 67.600 43.600 68.400 ;
        RECT 38.200 66.200 41.800 66.600 ;
        RECT 42.800 66.200 43.400 67.600 ;
        RECT 46.000 66.200 46.800 69.700 ;
        RECT 38.000 66.000 42.000 66.200 ;
        RECT 38.000 62.200 38.800 66.000 ;
        RECT 41.200 62.200 42.000 66.000 ;
        RECT 42.800 62.200 43.600 66.200 ;
        RECT 45.000 65.600 46.800 66.200 ;
        RECT 50.800 70.300 51.600 79.800 ;
        RECT 55.000 72.400 55.800 79.800 ;
        RECT 56.400 73.600 57.200 74.400 ;
        RECT 56.600 72.400 57.200 73.600 ;
        RECT 55.000 71.800 56.000 72.400 ;
        RECT 56.600 71.800 58.000 72.400 ;
        RECT 54.000 70.300 54.800 70.400 ;
        RECT 50.800 69.700 54.800 70.300 ;
        RECT 45.000 62.200 45.800 65.600 ;
        RECT 50.800 62.200 51.600 69.700 ;
        RECT 54.000 68.800 54.800 69.700 ;
        RECT 55.400 68.400 56.000 71.800 ;
        RECT 57.200 71.600 58.000 71.800 ;
        RECT 60.400 70.300 61.200 79.800 ;
        RECT 64.600 72.400 65.400 79.800 ;
        RECT 66.000 73.600 66.800 74.400 ;
        RECT 66.200 72.400 66.800 73.600 ;
        RECT 68.400 72.400 69.200 79.800 ;
        RECT 64.600 71.800 65.600 72.400 ;
        RECT 66.200 71.800 67.600 72.400 ;
        RECT 68.400 71.800 70.600 72.400 ;
        RECT 63.600 70.300 64.400 70.400 ;
        RECT 60.400 69.700 64.400 70.300 ;
        RECT 55.400 68.300 58.000 68.400 ;
        RECT 58.800 68.300 59.600 68.400 ;
        RECT 55.400 67.700 59.600 68.300 ;
        RECT 55.400 67.600 58.000 67.700 ;
        RECT 58.800 67.600 59.600 67.700 ;
        RECT 52.600 66.200 56.200 66.600 ;
        RECT 57.200 66.200 57.800 67.600 ;
        RECT 52.400 66.000 56.400 66.200 ;
        RECT 52.400 62.200 53.200 66.000 ;
        RECT 55.600 62.200 56.400 66.000 ;
        RECT 57.200 62.200 58.000 66.200 ;
        RECT 58.800 64.800 59.600 66.400 ;
        RECT 60.400 62.200 61.200 69.700 ;
        RECT 63.600 68.800 64.400 69.700 ;
        RECT 65.000 70.300 65.600 71.800 ;
        RECT 66.800 71.600 67.600 71.800 ;
        RECT 70.000 71.200 70.600 71.800 ;
        RECT 70.000 70.400 71.200 71.200 ;
        RECT 68.400 70.300 69.200 70.400 ;
        RECT 65.000 69.700 69.200 70.300 ;
        RECT 65.000 68.400 65.600 69.700 ;
        RECT 68.400 68.800 69.200 69.700 ;
        RECT 65.000 67.600 67.600 68.400 ;
        RECT 62.200 66.200 65.800 66.600 ;
        RECT 66.800 66.200 67.400 67.600 ;
        RECT 70.000 67.400 70.600 70.400 ;
        RECT 68.400 66.800 70.600 67.400 ;
        RECT 78.000 66.800 78.800 68.400 ;
        RECT 62.000 66.000 66.000 66.200 ;
        RECT 62.000 62.200 62.800 66.000 ;
        RECT 65.200 62.200 66.000 66.000 ;
        RECT 66.800 62.200 67.600 66.200 ;
        RECT 68.400 62.200 69.200 66.800 ;
        RECT 79.600 66.200 80.400 79.800 ;
        RECT 84.400 70.300 85.200 79.800 ;
        RECT 88.600 72.400 89.400 79.800 ;
        RECT 90.000 73.600 90.800 74.400 ;
        RECT 90.200 72.400 90.800 73.600 ;
        RECT 88.600 71.800 89.600 72.400 ;
        RECT 90.200 71.800 91.600 72.400 ;
        RECT 87.600 70.300 88.400 70.400 ;
        RECT 84.400 69.700 88.400 70.300 ;
        RECT 79.600 65.600 81.400 66.200 ;
        RECT 80.600 64.400 81.400 65.600 ;
        RECT 82.800 64.800 83.600 66.400 ;
        RECT 79.600 63.600 81.400 64.400 ;
        RECT 80.600 62.200 81.400 63.600 ;
        RECT 84.400 62.200 85.200 69.700 ;
        RECT 87.600 68.800 88.400 69.700 ;
        RECT 89.000 68.400 89.600 71.800 ;
        RECT 90.800 71.600 91.600 71.800 ;
        RECT 89.000 68.300 91.600 68.400 ;
        RECT 92.400 68.300 93.200 68.400 ;
        RECT 89.000 67.700 93.200 68.300 ;
        RECT 89.000 67.600 91.600 67.700 ;
        RECT 92.400 67.600 93.200 67.700 ;
        RECT 86.200 66.200 89.800 66.600 ;
        RECT 90.800 66.200 91.400 67.600 ;
        RECT 94.000 66.200 94.800 79.800 ;
        RECT 98.800 70.300 99.600 79.800 ;
        RECT 101.200 73.600 102.000 74.400 ;
        RECT 101.200 72.400 101.800 73.600 ;
        RECT 102.600 72.400 103.400 79.800 ;
        RECT 100.400 71.800 101.800 72.400 ;
        RECT 102.400 71.800 103.400 72.400 ;
        RECT 100.400 71.600 101.200 71.800 ;
        RECT 100.400 70.300 101.200 70.400 ;
        RECT 98.800 69.700 101.200 70.300 ;
        RECT 95.600 68.300 96.400 68.400 ;
        RECT 95.600 67.700 97.900 68.300 ;
        RECT 95.600 66.800 96.400 67.700 ;
        RECT 97.300 66.400 97.900 67.700 ;
        RECT 86.000 66.000 90.000 66.200 ;
        RECT 86.000 62.200 86.800 66.000 ;
        RECT 89.200 62.200 90.000 66.000 ;
        RECT 90.800 62.200 91.600 66.200 ;
        RECT 93.000 65.600 94.800 66.200 ;
        RECT 93.000 64.400 93.800 65.600 ;
        RECT 97.200 64.800 98.000 66.400 ;
        RECT 92.400 63.600 93.800 64.400 ;
        RECT 93.000 62.200 93.800 63.600 ;
        RECT 98.800 62.200 99.600 69.700 ;
        RECT 100.400 69.600 101.200 69.700 ;
        RECT 102.400 68.400 103.000 71.800 ;
        RECT 103.600 68.800 104.400 70.400 ;
        RECT 100.400 67.600 103.000 68.400 ;
        RECT 100.600 66.200 101.200 67.600 ;
        RECT 102.200 66.200 105.800 66.600 ;
        RECT 100.400 62.200 101.200 66.200 ;
        RECT 102.000 66.000 106.000 66.200 ;
        RECT 102.000 62.200 102.800 66.000 ;
        RECT 105.200 62.200 106.000 66.000 ;
        RECT 3.800 58.400 4.600 59.800 ;
        RECT 2.800 57.600 4.600 58.400 ;
        RECT 3.800 56.400 4.600 57.600 ;
        RECT 2.800 55.800 4.600 56.400 ;
        RECT 2.800 42.200 3.600 55.800 ;
        RECT 7.600 42.200 8.400 59.800 ;
        RECT 9.800 56.400 10.600 59.800 ;
        RECT 9.800 55.800 11.600 56.400 ;
        RECT 10.800 42.200 11.600 55.800 ;
        RECT 14.000 55.600 14.800 57.200 ;
        RECT 12.400 54.300 13.200 55.200 ;
        RECT 14.100 54.300 14.700 55.600 ;
        RECT 12.400 53.700 14.700 54.300 ;
        RECT 12.400 53.600 13.200 53.700 ;
        RECT 15.600 52.300 16.400 59.800 ;
        RECT 17.200 56.000 18.000 59.800 ;
        RECT 20.400 56.000 21.200 59.800 ;
        RECT 17.200 55.800 21.200 56.000 ;
        RECT 22.000 55.800 22.800 59.800 ;
        RECT 24.200 56.400 25.000 59.800 ;
        RECT 24.200 55.800 26.000 56.400 ;
        RECT 33.200 56.000 34.000 59.800 ;
        RECT 36.400 56.000 37.200 59.800 ;
        RECT 33.200 55.800 37.200 56.000 ;
        RECT 17.400 55.400 21.000 55.800 ;
        RECT 22.000 54.400 22.600 55.800 ;
        RECT 20.200 53.600 22.800 54.400 ;
        RECT 18.800 52.300 19.600 53.200 ;
        RECT 15.600 51.700 19.600 52.300 ;
        RECT 15.600 42.200 16.400 51.700 ;
        RECT 18.800 51.600 19.600 51.700 ;
        RECT 20.200 50.200 20.800 53.600 ;
        RECT 25.200 52.300 26.000 55.800 ;
        RECT 33.400 55.400 37.000 55.800 ;
        RECT 38.000 55.600 38.800 59.800 ;
        RECT 40.200 56.400 41.000 59.800 ;
        RECT 40.200 55.800 42.000 56.400 ;
        RECT 26.800 53.600 27.600 55.200 ;
        RECT 38.000 54.400 38.600 55.600 ;
        RECT 36.200 53.600 38.800 54.400 ;
        RECT 22.100 51.700 26.000 52.300 ;
        RECT 22.100 50.400 22.700 51.700 ;
        RECT 22.000 50.200 22.800 50.400 ;
        RECT 19.800 49.600 20.800 50.200 ;
        RECT 21.400 49.600 22.800 50.200 ;
        RECT 19.800 42.200 20.600 49.600 ;
        RECT 21.400 48.400 22.000 49.600 ;
        RECT 21.200 47.600 22.000 48.400 ;
        RECT 25.200 42.200 26.000 51.700 ;
        RECT 30.000 52.300 30.800 52.400 ;
        RECT 34.800 52.300 35.600 53.200 ;
        RECT 30.000 51.700 35.600 52.300 ;
        RECT 30.000 51.600 30.800 51.700 ;
        RECT 34.800 51.600 35.600 51.700 ;
        RECT 36.200 50.200 36.800 53.600 ;
        RECT 41.200 52.300 42.000 55.800 ;
        RECT 44.400 55.600 45.200 57.200 ;
        RECT 38.100 51.700 42.000 52.300 ;
        RECT 38.100 50.400 38.700 51.700 ;
        RECT 38.000 50.200 38.800 50.400 ;
        RECT 35.800 49.600 36.800 50.200 ;
        RECT 37.400 49.600 38.800 50.200 ;
        RECT 35.800 42.200 36.600 49.600 ;
        RECT 37.400 48.400 38.000 49.600 ;
        RECT 37.200 47.600 38.000 48.400 ;
        RECT 41.200 42.200 42.000 51.700 ;
        RECT 46.000 50.300 46.800 59.800 ;
        RECT 50.200 58.400 51.000 59.800 ;
        RECT 50.200 57.600 51.600 58.400 ;
        RECT 50.200 56.400 51.000 57.600 ;
        RECT 49.200 55.800 51.000 56.400 ;
        RECT 52.400 56.000 53.200 59.800 ;
        RECT 55.600 56.000 56.400 59.800 ;
        RECT 52.400 55.800 56.400 56.000 ;
        RECT 57.200 55.800 58.000 59.800 ;
        RECT 59.400 56.400 60.200 59.800 ;
        RECT 66.200 58.400 67.000 59.800 ;
        RECT 66.200 57.600 67.600 58.400 ;
        RECT 66.200 56.400 67.000 57.600 ;
        RECT 59.400 55.800 61.200 56.400 ;
        RECT 47.600 50.300 48.400 50.400 ;
        RECT 46.000 49.700 48.400 50.300 ;
        RECT 46.000 42.200 46.800 49.700 ;
        RECT 47.600 49.600 48.400 49.700 ;
        RECT 49.200 42.200 50.000 55.800 ;
        RECT 52.600 55.400 56.200 55.800 ;
        RECT 57.200 54.400 57.800 55.800 ;
        RECT 55.400 54.300 58.000 54.400 ;
        RECT 58.800 54.300 59.600 54.400 ;
        RECT 55.400 53.700 59.600 54.300 ;
        RECT 55.400 53.600 58.000 53.700 ;
        RECT 58.800 53.600 59.600 53.700 ;
        RECT 54.000 51.600 54.800 53.200 ;
        RECT 55.400 50.200 56.000 53.600 ;
        RECT 60.400 52.300 61.200 55.800 ;
        RECT 65.200 55.800 67.000 56.400 ;
        RECT 62.000 53.600 62.800 55.200 ;
        RECT 63.600 53.600 64.400 55.200 ;
        RECT 57.300 51.700 61.200 52.300 ;
        RECT 57.300 50.400 57.900 51.700 ;
        RECT 57.200 50.200 58.000 50.400 ;
        RECT 55.000 49.600 56.000 50.200 ;
        RECT 56.600 49.600 58.000 50.200 ;
        RECT 55.000 42.200 55.800 49.600 ;
        RECT 56.600 48.400 57.200 49.600 ;
        RECT 56.400 47.600 57.200 48.400 ;
        RECT 60.400 42.200 61.200 51.700 ;
        RECT 65.200 42.200 66.000 55.800 ;
        RECT 68.400 55.600 69.200 57.200 ;
        RECT 70.000 42.200 70.800 59.800 ;
        RECT 71.600 55.600 72.400 57.200 ;
        RECT 73.200 52.300 74.000 59.800 ;
        RECT 79.600 55.800 80.400 59.800 ;
        RECT 81.200 56.000 82.000 59.800 ;
        RECT 84.400 56.000 85.200 59.800 ;
        RECT 81.200 55.800 85.200 56.000 ;
        RECT 86.600 58.400 87.400 59.800 ;
        RECT 93.400 58.400 94.200 59.800 ;
        RECT 86.600 57.600 88.400 58.400 ;
        RECT 93.400 57.600 94.800 58.400 ;
        RECT 86.600 56.400 87.400 57.600 ;
        RECT 93.400 56.400 94.200 57.600 ;
        RECT 86.600 55.800 88.400 56.400 ;
        RECT 79.800 54.400 80.400 55.800 ;
        RECT 81.400 55.400 85.000 55.800 ;
        RECT 79.600 53.600 82.200 54.400 ;
        RECT 78.000 52.300 78.800 52.400 ;
        RECT 73.200 51.700 78.800 52.300 ;
        RECT 73.200 42.200 74.000 51.700 ;
        RECT 78.000 51.600 78.800 51.700 ;
        RECT 79.600 50.200 80.400 50.400 ;
        RECT 81.600 50.200 82.200 53.600 ;
        RECT 82.800 51.600 83.600 53.200 ;
        RECT 79.600 49.600 81.000 50.200 ;
        RECT 81.600 49.600 82.600 50.200 ;
        RECT 80.400 48.400 81.000 49.600 ;
        RECT 80.400 47.600 81.200 48.400 ;
        RECT 81.800 44.400 82.600 49.600 ;
        RECT 81.800 43.600 83.600 44.400 ;
        RECT 81.800 42.200 82.600 43.600 ;
        RECT 87.600 42.200 88.400 55.800 ;
        RECT 92.400 55.800 94.200 56.400 ;
        RECT 95.600 55.800 96.400 59.800 ;
        RECT 97.200 56.000 98.000 59.800 ;
        RECT 100.400 56.000 101.200 59.800 ;
        RECT 97.200 55.800 101.200 56.000 ;
        RECT 92.400 42.200 93.200 55.800 ;
        RECT 95.800 54.400 96.400 55.800 ;
        RECT 97.400 55.400 101.000 55.800 ;
        RECT 102.000 55.200 102.800 59.800 ;
        RECT 102.000 54.600 104.200 55.200 ;
        RECT 95.600 53.600 98.200 54.400 ;
        RECT 97.600 52.400 98.200 53.600 ;
        RECT 97.200 51.600 98.200 52.400 ;
        RECT 98.800 51.600 99.600 53.200 ;
        RECT 100.400 52.300 101.200 52.400 ;
        RECT 102.000 52.300 102.800 53.200 ;
        RECT 100.400 51.700 102.800 52.300 ;
        RECT 100.400 51.600 101.200 51.700 ;
        RECT 102.000 51.600 102.800 51.700 ;
        RECT 103.600 51.600 104.200 54.600 ;
        RECT 95.600 50.200 96.400 50.400 ;
        RECT 97.600 50.200 98.200 51.600 ;
        RECT 103.600 50.800 104.800 51.600 ;
        RECT 103.600 50.200 104.200 50.800 ;
        RECT 95.600 49.600 97.000 50.200 ;
        RECT 97.600 49.600 98.600 50.200 ;
        RECT 96.400 48.400 97.000 49.600 ;
        RECT 96.400 47.600 97.200 48.400 ;
        RECT 97.800 42.200 98.600 49.600 ;
        RECT 102.000 49.600 104.200 50.200 ;
        RECT 102.000 42.200 102.800 49.600 ;
        RECT 2.800 22.200 3.600 39.800 ;
        RECT 7.600 32.400 8.400 39.800 ;
        RECT 10.000 33.600 10.800 34.400 ;
        RECT 10.000 32.400 10.600 33.600 ;
        RECT 11.400 32.400 12.200 39.800 ;
        RECT 6.200 31.800 8.400 32.400 ;
        RECT 9.200 31.800 10.600 32.400 ;
        RECT 11.200 31.800 12.200 32.400 ;
        RECT 6.200 31.200 6.800 31.800 ;
        RECT 9.200 31.600 10.000 31.800 ;
        RECT 5.600 30.400 6.800 31.200 ;
        RECT 6.200 27.400 6.800 30.400 ;
        RECT 7.600 30.300 8.400 30.400 ;
        RECT 11.200 30.300 11.800 31.800 ;
        RECT 7.600 29.700 11.800 30.300 ;
        RECT 7.600 28.800 8.400 29.700 ;
        RECT 11.200 28.400 11.800 29.700 ;
        RECT 12.400 30.300 13.200 30.400 ;
        RECT 15.600 30.300 16.400 39.800 ;
        RECT 12.400 29.700 16.400 30.300 ;
        RECT 12.400 28.800 13.200 29.700 ;
        RECT 9.200 27.600 11.800 28.400 ;
        RECT 6.200 26.800 8.400 27.400 ;
        RECT 7.600 22.200 8.400 26.800 ;
        RECT 9.400 26.200 10.000 27.600 ;
        RECT 11.000 26.200 14.600 26.600 ;
        RECT 9.200 22.200 10.000 26.200 ;
        RECT 10.800 26.000 14.800 26.200 ;
        RECT 10.800 22.200 11.600 26.000 ;
        RECT 14.000 22.200 14.800 26.000 ;
        RECT 15.600 22.200 16.400 29.700 ;
        RECT 17.200 24.800 18.000 26.400 ;
        RECT 20.400 26.200 21.200 39.800 ;
        RECT 31.000 32.400 31.800 39.800 ;
        RECT 32.400 33.600 33.200 34.400 ;
        RECT 32.600 32.400 33.200 33.600 ;
        RECT 31.000 31.800 32.000 32.400 ;
        RECT 32.600 31.800 34.000 32.400 ;
        RECT 30.000 28.800 30.800 30.400 ;
        RECT 31.400 28.400 32.000 31.800 ;
        RECT 33.200 31.600 34.000 31.800 ;
        RECT 36.400 30.300 37.200 39.800 ;
        RECT 40.600 38.400 41.400 39.800 ;
        RECT 39.600 37.600 41.400 38.400 ;
        RECT 40.600 32.400 41.400 37.600 ;
        RECT 42.000 33.600 42.800 34.400 ;
        RECT 42.200 32.400 42.800 33.600 ;
        RECT 40.600 31.800 41.600 32.400 ;
        RECT 42.200 31.800 43.600 32.400 ;
        RECT 39.600 30.300 40.400 30.400 ;
        RECT 36.400 29.700 40.400 30.300 ;
        RECT 22.000 28.300 22.800 28.400 ;
        RECT 26.800 28.300 27.600 28.400 ;
        RECT 22.000 27.700 27.600 28.300 ;
        RECT 22.000 26.800 22.800 27.700 ;
        RECT 26.800 27.600 27.600 27.700 ;
        RECT 31.400 27.600 34.000 28.400 ;
        RECT 28.600 26.200 32.200 26.600 ;
        RECT 33.200 26.300 33.800 27.600 ;
        RECT 34.800 26.300 35.600 26.400 ;
        RECT 19.400 25.600 21.200 26.200 ;
        RECT 28.400 26.000 32.400 26.200 ;
        RECT 19.400 24.400 20.200 25.600 ;
        RECT 18.800 23.600 20.200 24.400 ;
        RECT 19.400 22.200 20.200 23.600 ;
        RECT 28.400 22.200 29.200 26.000 ;
        RECT 31.600 22.200 32.400 26.000 ;
        RECT 33.200 25.700 35.600 26.300 ;
        RECT 33.200 22.200 34.000 25.700 ;
        RECT 34.800 24.800 35.600 25.700 ;
        RECT 36.400 22.200 37.200 29.700 ;
        RECT 39.600 28.800 40.400 29.700 ;
        RECT 41.000 28.400 41.600 31.800 ;
        RECT 42.800 31.600 43.600 31.800 ;
        RECT 42.900 30.300 43.500 31.600 ;
        RECT 44.400 30.300 45.200 30.400 ;
        RECT 42.900 29.700 45.200 30.300 ;
        RECT 44.400 29.600 45.200 29.700 ;
        RECT 41.000 27.600 43.600 28.400 ;
        RECT 38.200 26.200 41.800 26.600 ;
        RECT 42.800 26.200 43.400 27.600 ;
        RECT 46.000 26.200 46.800 39.800 ;
        RECT 38.000 26.000 42.000 26.200 ;
        RECT 38.000 22.200 38.800 26.000 ;
        RECT 41.200 22.200 42.000 26.000 ;
        RECT 42.800 22.200 43.600 26.200 ;
        RECT 45.000 25.600 46.800 26.200 ;
        RECT 50.800 26.200 51.600 39.800 ;
        RECT 55.600 30.300 56.400 39.800 ;
        RECT 59.800 32.400 60.600 39.800 ;
        RECT 61.200 33.600 62.000 34.400 ;
        RECT 61.400 32.400 62.000 33.600 ;
        RECT 59.800 31.800 60.800 32.400 ;
        RECT 61.400 31.800 62.800 32.400 ;
        RECT 58.800 30.300 59.600 30.400 ;
        RECT 55.600 29.700 59.600 30.300 ;
        RECT 50.800 25.600 52.600 26.200 ;
        RECT 45.000 24.400 45.800 25.600 ;
        RECT 45.000 23.600 46.800 24.400 ;
        RECT 45.000 22.200 45.800 23.600 ;
        RECT 51.800 22.200 52.600 25.600 ;
        RECT 54.000 24.800 54.800 26.400 ;
        RECT 55.600 22.200 56.400 29.700 ;
        RECT 58.800 28.800 59.600 29.700 ;
        RECT 60.200 28.400 60.800 31.800 ;
        RECT 62.000 31.600 62.800 31.800 ;
        RECT 62.100 30.300 62.700 31.600 ;
        RECT 65.200 30.300 66.000 39.800 ;
        RECT 62.100 29.700 66.000 30.300 ;
        RECT 60.200 28.300 62.800 28.400 ;
        RECT 63.600 28.300 64.400 28.400 ;
        RECT 60.200 27.700 64.400 28.300 ;
        RECT 60.200 27.600 62.800 27.700 ;
        RECT 63.600 27.600 64.400 27.700 ;
        RECT 57.400 26.200 61.000 26.600 ;
        RECT 62.000 26.200 62.600 27.600 ;
        RECT 65.200 26.200 66.000 29.700 ;
        RECT 68.400 26.800 69.200 28.400 ;
        RECT 57.200 26.000 61.200 26.200 ;
        RECT 57.200 22.200 58.000 26.000 ;
        RECT 60.400 22.200 61.200 26.000 ;
        RECT 62.000 22.200 62.800 26.200 ;
        RECT 64.200 25.600 66.000 26.200 ;
        RECT 70.000 26.200 70.800 39.800 ;
        RECT 79.600 30.300 80.400 39.800 ;
        RECT 83.800 32.400 84.600 39.800 ;
        RECT 85.200 33.600 86.000 34.400 ;
        RECT 85.400 32.400 86.000 33.600 ;
        RECT 83.800 31.800 84.800 32.400 ;
        RECT 85.400 31.800 86.800 32.400 ;
        RECT 82.800 30.300 83.600 30.400 ;
        RECT 79.600 29.700 83.600 30.300 ;
        RECT 70.000 25.600 71.800 26.200 ;
        RECT 64.200 22.200 65.000 25.600 ;
        RECT 71.000 24.400 71.800 25.600 ;
        RECT 78.000 24.800 78.800 26.400 ;
        RECT 70.000 23.600 71.800 24.400 ;
        RECT 71.000 22.200 71.800 23.600 ;
        RECT 79.600 22.200 80.400 29.700 ;
        RECT 82.800 28.800 83.600 29.700 ;
        RECT 84.200 28.400 84.800 31.800 ;
        RECT 86.000 31.600 86.800 31.800 ;
        RECT 84.200 27.600 86.800 28.400 ;
        RECT 81.400 26.200 85.000 26.600 ;
        RECT 86.000 26.200 86.600 27.600 ;
        RECT 87.600 26.800 88.400 28.400 ;
        RECT 89.200 26.200 90.000 39.800 ;
        RECT 92.400 26.800 93.200 28.400 ;
        RECT 94.000 26.200 94.800 39.800 ;
        RECT 97.200 32.400 98.000 39.800 ;
        RECT 102.000 32.400 102.800 39.800 ;
        RECT 97.200 31.800 99.400 32.400 ;
        RECT 102.000 31.800 104.200 32.400 ;
        RECT 98.800 31.200 99.400 31.800 ;
        RECT 103.600 31.200 104.200 31.800 ;
        RECT 98.800 30.400 100.000 31.200 ;
        RECT 103.600 30.400 104.800 31.200 ;
        RECT 97.200 28.800 98.000 30.400 ;
        RECT 98.800 27.400 99.400 30.400 ;
        RECT 102.000 28.800 102.800 30.400 ;
        RECT 103.600 27.400 104.200 30.400 ;
        RECT 97.200 26.800 99.400 27.400 ;
        RECT 102.000 26.800 104.200 27.400 ;
        RECT 81.200 26.000 85.200 26.200 ;
        RECT 81.200 22.200 82.000 26.000 ;
        RECT 84.400 22.200 85.200 26.000 ;
        RECT 86.000 22.200 86.800 26.200 ;
        RECT 89.200 25.600 91.000 26.200 ;
        RECT 94.000 25.600 95.800 26.200 ;
        RECT 90.200 24.400 91.000 25.600 ;
        RECT 90.200 23.600 91.600 24.400 ;
        RECT 90.200 22.200 91.000 23.600 ;
        RECT 95.000 22.200 95.800 25.600 ;
        RECT 97.200 22.200 98.000 26.800 ;
        RECT 102.000 22.200 102.800 26.800 ;
        RECT 2.800 12.300 3.600 19.800 ;
        RECT 4.400 16.000 5.200 19.800 ;
        RECT 7.600 16.000 8.400 19.800 ;
        RECT 4.400 15.800 8.400 16.000 ;
        RECT 9.200 16.300 10.000 19.800 ;
        RECT 10.800 16.300 11.600 17.200 ;
        RECT 4.600 15.400 8.200 15.800 ;
        RECT 9.200 15.700 11.600 16.300 ;
        RECT 9.200 14.400 9.800 15.700 ;
        RECT 10.800 15.600 11.600 15.700 ;
        RECT 7.400 13.600 10.000 14.400 ;
        RECT 6.000 12.300 6.800 13.200 ;
        RECT 2.800 11.700 6.800 12.300 ;
        RECT 2.800 2.200 3.600 11.700 ;
        RECT 6.000 11.600 6.800 11.700 ;
        RECT 7.400 10.200 8.000 13.600 ;
        RECT 12.400 12.300 13.200 19.800 ;
        RECT 14.000 16.000 14.800 19.800 ;
        RECT 17.200 16.000 18.000 19.800 ;
        RECT 14.000 15.800 18.000 16.000 ;
        RECT 18.800 15.800 19.600 19.800 ;
        RECT 21.000 16.400 21.800 19.800 ;
        RECT 21.000 15.800 22.800 16.400 ;
        RECT 14.200 15.400 17.800 15.800 ;
        RECT 18.800 14.400 19.400 15.800 ;
        RECT 17.000 13.600 19.600 14.400 ;
        RECT 15.600 12.300 16.400 13.200 ;
        RECT 12.400 11.700 16.400 12.300 ;
        RECT 9.200 10.200 10.000 10.400 ;
        RECT 7.000 9.600 8.000 10.200 ;
        RECT 8.600 9.600 10.000 10.200 ;
        RECT 7.000 2.200 7.800 9.600 ;
        RECT 8.600 8.400 9.200 9.600 ;
        RECT 8.400 7.600 9.200 8.400 ;
        RECT 12.400 2.200 13.200 11.700 ;
        RECT 15.600 11.600 16.400 11.700 ;
        RECT 17.000 10.200 17.600 13.600 ;
        RECT 18.800 10.200 19.600 10.400 ;
        RECT 16.600 9.600 17.600 10.200 ;
        RECT 18.200 9.600 19.600 10.200 ;
        RECT 16.600 2.200 17.400 9.600 ;
        RECT 18.200 8.400 18.800 9.600 ;
        RECT 18.000 7.600 18.800 8.400 ;
        RECT 22.000 2.200 22.800 15.800 ;
        RECT 31.600 2.200 32.400 19.800 ;
        RECT 33.800 18.400 34.600 19.800 ;
        RECT 33.200 17.600 34.600 18.400 ;
        RECT 33.800 16.400 34.600 17.600 ;
        RECT 33.800 15.800 35.600 16.400 ;
        RECT 38.000 16.000 38.800 19.800 ;
        RECT 41.200 16.000 42.000 19.800 ;
        RECT 38.000 15.800 42.000 16.000 ;
        RECT 34.800 2.200 35.600 15.800 ;
        RECT 38.200 15.400 41.800 15.800 ;
        RECT 42.800 15.600 43.600 19.800 ;
        RECT 45.000 18.400 45.800 19.800 ;
        RECT 44.400 17.600 45.800 18.400 ;
        RECT 45.000 16.400 45.800 17.600 ;
        RECT 45.000 15.800 46.800 16.400 ;
        RECT 42.800 14.400 43.400 15.600 ;
        RECT 41.000 13.600 43.600 14.400 ;
        RECT 39.600 11.600 40.400 13.200 ;
        RECT 41.000 10.200 41.600 13.600 ;
        RECT 42.800 10.200 43.600 10.400 ;
        RECT 40.600 9.600 41.600 10.200 ;
        RECT 42.200 9.600 43.600 10.200 ;
        RECT 40.600 2.200 41.400 9.600 ;
        RECT 42.200 8.400 42.800 9.600 ;
        RECT 42.000 7.600 42.800 8.400 ;
        RECT 46.000 2.200 46.800 15.800 ;
        RECT 47.600 13.600 48.400 15.200 ;
        RECT 50.800 12.300 51.600 19.800 ;
        RECT 52.400 16.000 53.200 19.800 ;
        RECT 55.600 16.000 56.400 19.800 ;
        RECT 52.400 15.800 56.400 16.000 ;
        RECT 57.200 15.800 58.000 19.800 ;
        RECT 61.400 16.400 62.200 19.800 ;
        RECT 60.400 15.800 62.200 16.400 ;
        RECT 52.600 15.400 56.200 15.800 ;
        RECT 57.200 14.400 57.800 15.800 ;
        RECT 55.400 14.300 58.000 14.400 ;
        RECT 58.800 14.300 59.600 15.200 ;
        RECT 55.400 13.700 59.600 14.300 ;
        RECT 55.400 13.600 58.000 13.700 ;
        RECT 58.800 13.600 59.600 13.700 ;
        RECT 54.000 12.300 54.800 13.200 ;
        RECT 50.800 11.700 54.800 12.300 ;
        RECT 50.800 2.200 51.600 11.700 ;
        RECT 54.000 11.600 54.800 11.700 ;
        RECT 55.400 10.200 56.000 13.600 ;
        RECT 57.200 10.200 58.000 10.400 ;
        RECT 55.000 9.600 56.000 10.200 ;
        RECT 56.600 9.600 58.000 10.200 ;
        RECT 55.000 2.200 55.800 9.600 ;
        RECT 56.600 8.400 57.200 9.600 ;
        RECT 56.400 7.600 57.200 8.400 ;
        RECT 60.400 2.200 61.200 15.800 ;
        RECT 63.600 15.600 64.400 17.200 ;
        RECT 65.200 2.200 66.000 19.800 ;
        RECT 66.800 15.800 67.600 19.800 ;
        RECT 68.400 16.000 69.200 19.800 ;
        RECT 71.600 16.000 72.400 19.800 ;
        RECT 68.400 15.800 72.400 16.000 ;
        RECT 78.000 15.800 78.800 19.800 ;
        RECT 79.600 16.000 80.400 19.800 ;
        RECT 82.800 16.000 83.600 19.800 ;
        RECT 79.600 15.800 83.600 16.000 ;
        RECT 67.000 14.400 67.600 15.800 ;
        RECT 68.600 15.400 72.200 15.800 ;
        RECT 78.200 14.400 78.800 15.800 ;
        RECT 79.800 15.400 83.400 15.800 ;
        RECT 66.800 13.600 69.400 14.400 ;
        RECT 78.000 13.600 80.600 14.400 ;
        RECT 66.800 10.200 67.600 10.400 ;
        RECT 68.800 10.200 69.400 13.600 ;
        RECT 70.000 11.600 70.800 13.200 ;
        RECT 80.000 12.400 80.600 13.600 ;
        RECT 79.600 11.600 80.600 12.400 ;
        RECT 81.200 12.300 82.000 13.200 ;
        RECT 84.400 12.300 85.200 19.800 ;
        RECT 86.000 15.600 86.800 17.200 ;
        RECT 87.600 15.200 88.400 19.800 ;
        RECT 92.400 15.600 93.200 17.200 ;
        RECT 87.600 14.600 89.800 15.200 ;
        RECT 81.200 11.700 85.200 12.300 ;
        RECT 81.200 11.600 82.000 11.700 ;
        RECT 78.000 10.200 78.800 10.400 ;
        RECT 80.000 10.200 80.600 11.600 ;
        RECT 66.800 9.600 68.200 10.200 ;
        RECT 68.800 9.600 69.800 10.200 ;
        RECT 78.000 9.600 79.400 10.200 ;
        RECT 80.000 9.600 81.000 10.200 ;
        RECT 67.600 8.400 68.200 9.600 ;
        RECT 67.600 7.600 68.400 8.400 ;
        RECT 69.000 2.200 69.800 9.600 ;
        RECT 78.800 8.400 79.400 9.600 ;
        RECT 78.800 7.600 79.600 8.400 ;
        RECT 80.200 2.200 81.000 9.600 ;
        RECT 84.400 2.200 85.200 11.700 ;
        RECT 86.000 12.300 86.800 12.400 ;
        RECT 87.600 12.300 88.400 13.200 ;
        RECT 86.000 11.700 88.400 12.300 ;
        RECT 86.000 11.600 86.800 11.700 ;
        RECT 87.600 11.600 88.400 11.700 ;
        RECT 89.200 11.600 89.800 14.600 ;
        RECT 89.200 10.800 90.400 11.600 ;
        RECT 89.200 10.200 89.800 10.800 ;
        RECT 87.600 9.600 89.800 10.200 ;
        RECT 87.600 2.200 88.400 9.600 ;
        RECT 94.000 2.200 94.800 19.800 ;
        RECT 95.600 15.800 96.400 19.800 ;
        RECT 97.200 16.000 98.000 19.800 ;
        RECT 100.400 16.000 101.200 19.800 ;
        RECT 97.200 15.800 101.200 16.000 ;
        RECT 95.800 14.400 96.400 15.800 ;
        RECT 97.400 15.400 101.000 15.800 ;
        RECT 102.000 15.200 102.800 19.800 ;
        RECT 102.000 14.600 104.200 15.200 ;
        RECT 95.600 13.600 98.200 14.400 ;
        RECT 97.600 12.400 98.200 13.600 ;
        RECT 97.200 11.600 98.200 12.400 ;
        RECT 98.800 11.600 99.600 13.200 ;
        RECT 100.400 12.300 101.200 12.400 ;
        RECT 102.000 12.300 102.800 13.200 ;
        RECT 100.400 11.700 102.800 12.300 ;
        RECT 100.400 11.600 101.200 11.700 ;
        RECT 102.000 11.600 102.800 11.700 ;
        RECT 103.600 11.600 104.200 14.600 ;
        RECT 95.600 10.200 96.400 10.400 ;
        RECT 97.600 10.200 98.200 11.600 ;
        RECT 103.600 10.800 104.800 11.600 ;
        RECT 103.600 10.200 104.200 10.800 ;
        RECT 95.600 9.600 97.000 10.200 ;
        RECT 97.600 9.600 98.600 10.200 ;
        RECT 96.400 8.400 97.000 9.600 ;
        RECT 96.400 7.600 97.200 8.400 ;
        RECT 97.800 2.200 98.600 9.600 ;
        RECT 102.000 9.600 104.200 10.200 ;
        RECT 102.000 2.200 102.800 9.600 ;
      LAYER via1 ;
        RECT 41.200 67.600 42.000 68.400 ;
        RECT 58.800 65.600 59.600 66.400 ;
        RECT 78.000 67.600 78.800 68.400 ;
        RECT 82.800 65.600 83.600 66.400 ;
        RECT 95.600 67.600 96.400 68.400 ;
        RECT 103.600 69.600 104.400 70.400 ;
        RECT 102.000 67.600 102.800 68.400 ;
        RECT 7.600 49.600 8.400 50.400 ;
        RECT 10.800 43.600 11.600 44.400 ;
        RECT 22.000 57.600 22.800 58.400 ;
        RECT 50.800 57.600 51.600 58.400 ;
        RECT 66.800 57.600 67.600 58.400 ;
        RECT 70.000 49.600 70.800 50.400 ;
        RECT 87.600 57.600 88.400 58.400 ;
        RECT 94.000 57.600 94.800 58.400 ;
        RECT 82.800 43.600 83.600 44.400 ;
        RECT 2.800 29.600 3.600 30.400 ;
        RECT 17.200 25.600 18.000 26.400 ;
        RECT 30.000 29.600 30.800 30.400 ;
        RECT 31.600 27.600 32.400 28.400 ;
        RECT 46.000 23.600 46.800 24.400 ;
        RECT 54.000 25.600 54.800 26.400 ;
        RECT 68.400 27.600 69.200 28.400 ;
        RECT 78.000 25.600 78.800 26.400 ;
        RECT 86.000 27.600 86.800 28.400 ;
        RECT 87.600 27.600 88.400 28.400 ;
        RECT 94.000 37.600 94.800 38.400 ;
        RECT 92.400 27.600 93.200 28.400 ;
        RECT 97.200 29.600 98.000 30.400 ;
        RECT 102.000 29.600 102.800 30.400 ;
        RECT 90.800 23.600 91.600 24.400 ;
        RECT 17.200 13.600 18.000 14.400 ;
        RECT 9.200 9.600 10.000 10.400 ;
        RECT 18.800 9.600 19.600 10.400 ;
        RECT 22.000 9.600 22.800 10.400 ;
        RECT 31.600 11.600 32.400 12.400 ;
        RECT 42.800 9.600 43.600 10.400 ;
        RECT 55.600 13.600 56.400 14.400 ;
        RECT 57.200 9.600 58.000 10.400 ;
        RECT 60.400 7.600 61.200 8.400 ;
        RECT 68.400 13.600 69.200 14.400 ;
        RECT 65.200 9.600 66.000 10.400 ;
        RECT 94.000 9.600 94.800 10.400 ;
      LAYER metal2 ;
        RECT 94.000 73.600 94.800 74.400 ;
        RECT 100.400 73.600 101.200 74.400 ;
        RECT 2.800 71.600 3.600 72.400 ;
        RECT 9.200 71.600 10.000 72.400 ;
        RECT 15.600 71.600 16.400 72.400 ;
        RECT 50.800 71.600 51.600 72.400 ;
        RECT 57.200 71.600 58.000 72.400 ;
        RECT 66.800 71.600 67.600 72.400 ;
        RECT 87.600 71.600 88.400 72.400 ;
        RECT 90.800 71.600 91.600 72.400 ;
        RECT 2.900 58.400 3.500 71.600 ;
        RECT 2.800 57.600 3.600 58.400 ;
        RECT 15.700 58.300 16.300 71.600 ;
        RECT 23.600 69.600 24.400 70.400 ;
        RECT 14.100 57.700 16.300 58.300 ;
        RECT 22.000 58.300 22.800 58.400 ;
        RECT 23.700 58.300 24.300 69.600 ;
        RECT 28.400 67.600 29.200 68.400 ;
        RECT 41.200 67.600 42.000 68.400 ;
        RECT 26.800 65.600 27.600 66.400 ;
        RECT 22.000 57.700 24.300 58.300 ;
        RECT 14.100 56.400 14.700 57.700 ;
        RECT 22.000 57.600 22.800 57.700 ;
        RECT 14.000 55.600 14.800 56.400 ;
        RECT 26.900 54.400 27.500 65.600 ;
        RECT 41.300 58.400 41.900 67.600 ;
        RECT 50.900 58.400 51.500 71.600 ;
        RECT 58.800 67.600 59.600 68.400 ;
        RECT 58.800 65.600 59.600 66.400 ;
        RECT 66.900 58.400 67.500 71.600 ;
        RECT 78.000 67.600 78.800 68.400 ;
        RECT 82.800 65.600 83.600 66.400 ;
        RECT 79.600 63.600 80.400 64.400 ;
        RECT 41.200 57.600 42.000 58.400 ;
        RECT 44.400 57.600 45.200 58.400 ;
        RECT 50.800 57.600 51.600 58.400 ;
        RECT 66.800 57.600 67.600 58.400 ;
        RECT 44.500 56.400 45.100 57.600 ;
        RECT 38.000 55.600 38.800 56.400 ;
        RECT 44.400 55.600 45.200 56.400 ;
        RECT 62.000 55.600 62.800 56.400 ;
        RECT 68.400 55.600 69.200 56.400 ;
        RECT 71.600 55.600 72.400 56.400 ;
        RECT 62.100 54.400 62.700 55.600 ;
        RECT 71.700 54.400 72.300 55.600 ;
        RECT 26.800 53.600 27.600 54.400 ;
        RECT 58.800 53.600 59.600 54.400 ;
        RECT 62.000 53.600 62.800 54.400 ;
        RECT 63.600 53.600 64.400 54.400 ;
        RECT 71.600 53.600 72.400 54.400 ;
        RECT 7.600 49.600 8.400 50.400 ;
        RECT 26.900 44.400 27.500 53.600 ;
        RECT 30.000 51.600 30.800 52.400 ;
        RECT 54.000 51.600 54.800 52.400 ;
        RECT 78.000 51.600 78.800 52.400 ;
        RECT 30.100 50.400 30.700 51.600 ;
        RECT 54.100 50.400 54.700 51.600 ;
        RECT 79.700 50.400 80.300 63.600 ;
        RECT 87.700 58.400 88.300 71.600 ;
        RECT 92.400 67.600 93.200 68.400 ;
        RECT 92.400 63.600 93.200 64.400 ;
        RECT 87.600 57.600 88.400 58.400 ;
        RECT 82.800 51.600 83.600 52.400 ;
        RECT 82.900 50.400 83.500 51.600 ;
        RECT 30.000 49.600 30.800 50.400 ;
        RECT 47.600 49.600 48.400 50.400 ;
        RECT 54.000 49.600 54.800 50.400 ;
        RECT 70.000 49.600 70.800 50.400 ;
        RECT 79.600 49.600 80.400 50.400 ;
        RECT 82.800 49.600 83.600 50.400 ;
        RECT 10.800 43.600 11.600 44.400 ;
        RECT 26.800 43.600 27.600 44.400 ;
        RECT 39.600 43.600 40.400 44.400 ;
        RECT 82.800 43.600 83.600 44.400 ;
        RECT 9.200 32.300 10.000 32.400 ;
        RECT 10.900 32.300 11.500 43.600 ;
        RECT 39.700 38.400 40.300 43.600 ;
        RECT 39.600 37.600 40.400 38.400 ;
        RECT 82.900 34.400 83.500 43.600 ;
        RECT 82.800 33.600 83.600 34.400 ;
        RECT 87.600 33.600 88.400 34.400 ;
        RECT 9.200 31.700 11.500 32.300 ;
        RECT 9.200 31.600 10.000 31.700 ;
        RECT 33.200 31.600 34.000 32.400 ;
        RECT 86.000 31.600 86.800 32.400 ;
        RECT 2.800 29.600 3.600 30.400 ;
        RECT 30.000 29.600 30.800 30.400 ;
        RECT 26.800 27.600 27.600 28.400 ;
        RECT 31.600 27.600 32.400 28.400 ;
        RECT 17.200 25.600 18.000 26.400 ;
        RECT 17.300 14.400 17.900 25.600 ;
        RECT 18.800 23.600 19.600 24.400 ;
        RECT 17.200 13.600 18.000 14.400 ;
        RECT 18.900 10.400 19.500 23.600 ;
        RECT 33.300 18.400 33.900 31.600 ;
        RECT 44.400 29.600 45.200 30.400 ;
        RECT 44.500 18.400 45.100 29.600 ;
        RECT 87.700 28.400 88.300 33.600 ;
        RECT 92.500 32.400 93.100 63.600 ;
        RECT 94.100 58.400 94.700 73.600 ;
        RECT 100.500 72.400 101.100 73.600 ;
        RECT 100.400 71.600 101.200 72.400 ;
        RECT 100.400 69.600 101.200 70.400 ;
        RECT 103.600 69.600 104.400 70.400 ;
        RECT 95.600 67.600 96.400 68.400 ;
        RECT 102.000 67.600 102.800 68.400 ;
        RECT 94.000 57.600 94.800 58.400 ;
        RECT 97.200 51.600 98.000 52.400 ;
        RECT 98.800 51.600 99.600 52.400 ;
        RECT 100.400 51.600 101.200 52.400 ;
        RECT 98.900 50.400 99.500 51.600 ;
        RECT 95.600 49.600 96.400 50.400 ;
        RECT 98.800 49.600 99.600 50.400 ;
        RECT 95.700 48.400 96.300 49.600 ;
        RECT 95.600 47.600 96.400 48.400 ;
        RECT 94.000 43.600 94.800 44.400 ;
        RECT 94.100 38.400 94.700 43.600 ;
        RECT 94.000 37.600 94.800 38.400 ;
        RECT 92.400 31.600 93.200 32.400 ;
        RECT 102.100 30.400 102.700 67.600 ;
        RECT 97.200 29.600 98.000 30.400 ;
        RECT 102.000 29.600 102.800 30.400 ;
        RECT 97.300 28.400 97.900 29.600 ;
        RECT 63.600 27.600 64.400 28.400 ;
        RECT 68.400 27.600 69.200 28.400 ;
        RECT 78.000 27.600 78.800 28.400 ;
        RECT 86.000 27.600 86.800 28.400 ;
        RECT 87.600 27.600 88.400 28.400 ;
        RECT 92.400 27.600 93.200 28.400 ;
        RECT 97.200 27.600 98.000 28.400 ;
        RECT 78.100 26.400 78.700 27.600 ;
        RECT 50.800 25.600 51.600 26.400 ;
        RECT 54.000 26.300 54.800 26.400 ;
        RECT 54.000 25.700 56.300 26.300 ;
        RECT 54.000 25.600 54.800 25.700 ;
        RECT 50.900 24.400 51.500 25.600 ;
        RECT 46.000 23.600 46.800 24.400 ;
        RECT 50.800 23.600 51.600 24.400 ;
        RECT 33.200 17.600 34.000 18.400 ;
        RECT 44.400 17.600 45.200 18.400 ;
        RECT 42.800 15.600 43.600 16.400 ;
        RECT 31.600 11.600 32.400 12.400 ;
        RECT 39.600 11.600 40.400 12.400 ;
        RECT 46.100 10.400 46.700 23.600 ;
        RECT 47.600 15.600 48.400 16.400 ;
        RECT 47.700 14.400 48.300 15.600 ;
        RECT 55.700 14.400 56.300 25.700 ;
        RECT 78.000 25.600 78.800 26.400 ;
        RECT 57.200 23.600 58.000 24.400 ;
        RECT 70.000 23.600 70.800 24.400 ;
        RECT 47.600 13.600 48.400 14.400 ;
        RECT 55.600 13.600 56.400 14.400 ;
        RECT 57.300 10.400 57.900 23.600 ;
        RECT 63.600 15.600 64.400 16.400 ;
        RECT 68.400 15.600 69.200 16.400 ;
        RECT 68.500 14.400 69.100 15.600 ;
        RECT 70.100 14.400 70.700 23.600 ;
        RECT 86.000 16.300 86.800 16.400 ;
        RECT 87.700 16.300 88.300 27.600 ;
        RECT 90.800 23.600 91.600 24.400 ;
        RECT 86.000 15.700 88.300 16.300 ;
        RECT 86.000 15.600 86.800 15.700 ;
        RECT 68.400 13.600 69.200 14.400 ;
        RECT 70.000 13.600 70.800 14.400 ;
        RECT 78.000 13.600 78.800 14.400 ;
        RECT 70.000 11.600 70.800 12.400 ;
        RECT 70.100 10.400 70.700 11.600 ;
        RECT 78.100 10.400 78.700 13.600 ;
        RECT 90.900 12.400 91.500 23.600 ;
        RECT 92.500 16.400 93.100 27.600 ;
        RECT 92.400 15.600 93.200 16.400 ;
        RECT 79.600 11.600 80.400 12.400 ;
        RECT 86.000 11.600 86.800 12.400 ;
        RECT 90.800 11.600 91.600 12.400 ;
        RECT 95.600 11.600 96.400 12.400 ;
        RECT 97.200 11.600 98.000 12.400 ;
        RECT 98.800 11.600 99.600 12.400 ;
        RECT 100.400 11.600 101.200 12.400 ;
        RECT 95.700 10.400 96.300 11.600 ;
        RECT 98.900 10.400 99.500 11.600 ;
        RECT 9.200 9.600 10.000 10.400 ;
        RECT 18.800 9.600 19.600 10.400 ;
        RECT 22.000 9.600 22.800 10.400 ;
        RECT 42.800 9.600 43.600 10.400 ;
        RECT 46.000 9.600 46.800 10.400 ;
        RECT 57.200 9.600 58.000 10.400 ;
        RECT 65.200 9.600 66.000 10.400 ;
        RECT 66.800 9.600 67.600 10.400 ;
        RECT 70.000 9.600 70.800 10.400 ;
        RECT 78.000 9.600 78.800 10.400 ;
        RECT 94.000 9.600 94.800 10.400 ;
        RECT 95.600 9.600 96.400 10.400 ;
        RECT 98.800 9.600 99.600 10.400 ;
        RECT 66.900 8.400 67.500 9.600 ;
        RECT 60.400 7.600 61.200 8.400 ;
        RECT 66.800 7.600 67.600 8.400 ;
      LAYER metal3 ;
        RECT 94.000 74.300 94.800 74.400 ;
        RECT 100.400 74.300 101.200 74.400 ;
        RECT 94.000 73.700 101.200 74.300 ;
        RECT 94.000 73.600 94.800 73.700 ;
        RECT 100.400 73.600 101.200 73.700 ;
        RECT 2.800 72.300 3.600 72.400 ;
        RECT 9.200 72.300 10.000 72.400 ;
        RECT 2.800 71.700 10.000 72.300 ;
        RECT 2.800 71.600 3.600 71.700 ;
        RECT 9.200 71.600 10.000 71.700 ;
        RECT 50.800 72.300 51.600 72.400 ;
        RECT 57.200 72.300 58.000 72.400 ;
        RECT 50.800 71.700 58.000 72.300 ;
        RECT 50.800 71.600 51.600 71.700 ;
        RECT 57.200 71.600 58.000 71.700 ;
        RECT 87.600 72.300 88.400 72.400 ;
        RECT 90.800 72.300 91.600 72.400 ;
        RECT 87.600 71.700 91.600 72.300 ;
        RECT 87.600 71.600 88.400 71.700 ;
        RECT 90.800 71.600 91.600 71.700 ;
        RECT 100.400 70.300 101.200 70.400 ;
        RECT 103.600 70.300 104.400 70.400 ;
        RECT 100.400 69.700 104.400 70.300 ;
        RECT 100.400 69.600 101.200 69.700 ;
        RECT 103.600 69.600 104.400 69.700 ;
        RECT 28.400 68.300 29.200 68.400 ;
        RECT 41.200 68.300 42.000 68.400 ;
        RECT 28.400 67.700 42.000 68.300 ;
        RECT 28.400 67.600 29.200 67.700 ;
        RECT 41.200 67.600 42.000 67.700 ;
        RECT 58.800 68.300 59.600 68.400 ;
        RECT 78.000 68.300 78.800 68.400 ;
        RECT 58.800 67.700 78.800 68.300 ;
        RECT 58.800 67.600 59.600 67.700 ;
        RECT 78.000 67.600 78.800 67.700 ;
        RECT 92.400 68.300 93.200 68.400 ;
        RECT 95.600 68.300 96.400 68.400 ;
        RECT 92.400 67.700 96.400 68.300 ;
        RECT 92.400 67.600 93.200 67.700 ;
        RECT 95.600 67.600 96.400 67.700 ;
        RECT 26.800 66.300 27.600 66.400 ;
        RECT 58.800 66.300 59.600 66.400 ;
        RECT 26.800 65.700 59.600 66.300 ;
        RECT 78.100 66.300 78.700 67.600 ;
        RECT 82.800 66.300 83.600 66.400 ;
        RECT 78.100 65.700 83.600 66.300 ;
        RECT 26.800 65.600 27.600 65.700 ;
        RECT 58.800 65.600 59.600 65.700 ;
        RECT 82.800 65.600 83.600 65.700 ;
        RECT 41.200 58.300 42.000 58.400 ;
        RECT 44.400 58.300 45.200 58.400 ;
        RECT 41.200 57.700 45.200 58.300 ;
        RECT 41.200 57.600 42.000 57.700 ;
        RECT 44.400 57.600 45.200 57.700 ;
        RECT 38.000 56.300 38.800 56.400 ;
        RECT 62.000 56.300 62.800 56.400 ;
        RECT 68.400 56.300 69.200 56.400 ;
        RECT 38.000 55.700 69.200 56.300 ;
        RECT 38.000 55.600 38.800 55.700 ;
        RECT 62.000 55.600 62.800 55.700 ;
        RECT 68.400 55.600 69.200 55.700 ;
        RECT 58.800 54.300 59.600 54.400 ;
        RECT 63.600 54.300 64.400 54.400 ;
        RECT 71.600 54.300 72.400 54.400 ;
        RECT 58.800 53.700 72.400 54.300 ;
        RECT 58.800 53.600 59.600 53.700 ;
        RECT 63.600 53.600 64.400 53.700 ;
        RECT 71.600 53.600 72.400 53.700 ;
        RECT 78.000 52.300 78.800 52.400 ;
        RECT 97.200 52.300 98.000 52.400 ;
        RECT 100.400 52.300 101.200 52.400 ;
        RECT 78.000 51.700 96.300 52.300 ;
        RECT 78.000 51.600 78.800 51.700 ;
        RECT 7.600 50.300 8.400 50.400 ;
        RECT 30.000 50.300 30.800 50.400 ;
        RECT 7.600 49.700 30.800 50.300 ;
        RECT 7.600 49.600 8.400 49.700 ;
        RECT 30.000 49.600 30.800 49.700 ;
        RECT 47.600 50.300 48.400 50.400 ;
        RECT 54.000 50.300 54.800 50.400 ;
        RECT 47.600 49.700 54.800 50.300 ;
        RECT 47.600 49.600 48.400 49.700 ;
        RECT 54.000 49.600 54.800 49.700 ;
        RECT 70.000 50.300 70.800 50.400 ;
        RECT 82.800 50.300 83.600 50.400 ;
        RECT 70.000 49.700 83.600 50.300 ;
        RECT 95.700 50.300 96.300 51.700 ;
        RECT 97.200 51.700 101.200 52.300 ;
        RECT 97.200 51.600 98.000 51.700 ;
        RECT 100.400 51.600 101.200 51.700 ;
        RECT 98.800 50.300 99.600 50.400 ;
        RECT 95.700 49.700 99.600 50.300 ;
        RECT 70.000 49.600 70.800 49.700 ;
        RECT 82.800 49.600 83.600 49.700 ;
        RECT 98.800 49.600 99.600 49.700 ;
        RECT 94.000 48.300 94.800 48.400 ;
        RECT 95.600 48.300 96.400 48.400 ;
        RECT 94.000 47.700 96.400 48.300 ;
        RECT 94.000 47.600 94.800 47.700 ;
        RECT 95.600 47.600 96.400 47.700 ;
        RECT 26.800 44.300 27.600 44.400 ;
        RECT 39.600 44.300 40.400 44.400 ;
        RECT 26.800 43.700 40.400 44.300 ;
        RECT 26.800 43.600 27.600 43.700 ;
        RECT 39.600 43.600 40.400 43.700 ;
        RECT 94.000 43.600 94.800 44.400 ;
        RECT 82.800 34.300 83.600 34.400 ;
        RECT 87.600 34.300 88.400 34.400 ;
        RECT 82.800 33.700 88.400 34.300 ;
        RECT 82.800 33.600 83.600 33.700 ;
        RECT 87.600 33.600 88.400 33.700 ;
        RECT 86.000 32.300 86.800 32.400 ;
        RECT 92.400 32.300 93.200 32.400 ;
        RECT 86.000 31.700 93.200 32.300 ;
        RECT 86.000 31.600 86.800 31.700 ;
        RECT 92.400 31.600 93.200 31.700 ;
        RECT 2.800 30.300 3.600 30.400 ;
        RECT 30.000 30.300 30.800 30.400 ;
        RECT 2.800 29.700 30.800 30.300 ;
        RECT 2.800 29.600 3.600 29.700 ;
        RECT 30.000 29.600 30.800 29.700 ;
        RECT 26.800 28.300 27.600 28.400 ;
        RECT 31.600 28.300 32.400 28.400 ;
        RECT 26.800 27.700 32.400 28.300 ;
        RECT 26.800 27.600 27.600 27.700 ;
        RECT 31.600 27.600 32.400 27.700 ;
        RECT 63.600 28.300 64.400 28.400 ;
        RECT 68.400 28.300 69.200 28.400 ;
        RECT 78.000 28.300 78.800 28.400 ;
        RECT 63.600 27.700 78.800 28.300 ;
        RECT 63.600 27.600 64.400 27.700 ;
        RECT 68.400 27.600 69.200 27.700 ;
        RECT 78.000 27.600 78.800 27.700 ;
        RECT 86.000 28.300 86.800 28.400 ;
        RECT 97.200 28.300 98.000 28.400 ;
        RECT 86.000 27.700 98.000 28.300 ;
        RECT 86.000 27.600 86.800 27.700 ;
        RECT 97.200 27.600 98.000 27.700 ;
        RECT 50.800 24.300 51.600 24.400 ;
        RECT 57.200 24.300 58.000 24.400 ;
        RECT 50.800 23.700 58.000 24.300 ;
        RECT 50.800 23.600 51.600 23.700 ;
        RECT 57.200 23.600 58.000 23.700 ;
        RECT 42.800 16.300 43.600 16.400 ;
        RECT 47.600 16.300 48.400 16.400 ;
        RECT 63.600 16.300 64.400 16.400 ;
        RECT 42.800 15.700 64.400 16.300 ;
        RECT 42.800 15.600 43.600 15.700 ;
        RECT 47.600 15.600 48.400 15.700 ;
        RECT 63.600 15.600 64.400 15.700 ;
        RECT 68.400 16.300 69.200 16.400 ;
        RECT 92.400 16.300 93.200 16.400 ;
        RECT 68.400 15.700 93.200 16.300 ;
        RECT 68.400 15.600 69.200 15.700 ;
        RECT 92.400 15.600 93.200 15.700 ;
        RECT 70.000 14.300 70.800 14.400 ;
        RECT 78.000 14.300 78.800 14.400 ;
        RECT 70.000 13.700 78.800 14.300 ;
        RECT 70.000 13.600 70.800 13.700 ;
        RECT 78.000 13.600 78.800 13.700 ;
        RECT 31.600 12.300 32.400 12.400 ;
        RECT 39.600 12.300 40.400 12.400 ;
        RECT 31.600 11.700 40.400 12.300 ;
        RECT 31.600 11.600 32.400 11.700 ;
        RECT 39.600 11.600 40.400 11.700 ;
        RECT 79.600 12.300 80.400 12.400 ;
        RECT 86.000 12.300 86.800 12.400 ;
        RECT 79.600 11.700 86.800 12.300 ;
        RECT 79.600 11.600 80.400 11.700 ;
        RECT 86.000 11.600 86.800 11.700 ;
        RECT 90.800 12.300 91.600 12.400 ;
        RECT 95.600 12.300 96.400 12.400 ;
        RECT 90.800 11.700 96.400 12.300 ;
        RECT 90.800 11.600 91.600 11.700 ;
        RECT 95.600 11.600 96.400 11.700 ;
        RECT 97.200 12.300 98.000 12.400 ;
        RECT 100.400 12.300 101.200 12.400 ;
        RECT 97.200 11.700 101.200 12.300 ;
        RECT 97.200 11.600 98.000 11.700 ;
        RECT 100.400 11.600 101.200 11.700 ;
        RECT 9.200 10.300 10.000 10.400 ;
        RECT 22.000 10.300 22.800 10.400 ;
        RECT 9.200 9.700 22.800 10.300 ;
        RECT 9.200 9.600 10.000 9.700 ;
        RECT 22.000 9.600 22.800 9.700 ;
        RECT 42.800 10.300 43.600 10.400 ;
        RECT 46.000 10.300 46.800 10.400 ;
        RECT 42.800 9.700 46.800 10.300 ;
        RECT 42.800 9.600 43.600 9.700 ;
        RECT 46.000 9.600 46.800 9.700 ;
        RECT 65.200 10.300 66.000 10.400 ;
        RECT 70.000 10.300 70.800 10.400 ;
        RECT 65.200 9.700 70.800 10.300 ;
        RECT 65.200 9.600 66.000 9.700 ;
        RECT 70.000 9.600 70.800 9.700 ;
        RECT 94.000 10.300 94.800 10.400 ;
        RECT 98.800 10.300 99.600 10.400 ;
        RECT 94.000 9.700 99.600 10.300 ;
        RECT 94.000 9.600 94.800 9.700 ;
        RECT 98.800 9.600 99.600 9.700 ;
        RECT 60.400 8.300 61.200 8.400 ;
        RECT 66.800 8.300 67.600 8.400 ;
        RECT 60.400 7.700 67.600 8.300 ;
        RECT 60.400 7.600 61.200 7.700 ;
        RECT 66.800 7.600 67.600 7.700 ;
      LAYER metal4 ;
        RECT 93.800 43.400 95.000 48.600 ;
  END
END barrel_shifter_8bit
END LIBRARY

